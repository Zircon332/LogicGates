<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-250.53,-402.064,261.95,-660.142</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>280.5,60.5</position>
<gparam>LABEL_TEXT Parallel and Serial Converter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>44,13</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>141.5,-41</position>
<gparam>LABEL_TEXT Color Storage</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>-228.5,-532</position>
<input>
<ID>IN_0</ID>459 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>46.5,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>775</ID>
<type>AA_LABEL</type>
<position>-221.5,-343</position>
<gparam>LABEL_TEXT Better Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-60,-300.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>50.5,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-235.5,-482.5</position>
<output>
<ID>OUT_0</ID>498 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>48.5,20</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>778</ID>
<type>BB_CLOCK</type>
<position>-234,-383</position>
<output>
<ID>CLK</ID>773 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-44,-21.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>779</ID>
<type>AA_AND2</type>
<position>-211,-381.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>773 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>32,19.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>780</ID>
<type>AA_REGISTER4</type>
<position>-212.5,-373.5</position>
<output>
<ID>OUT_0</ID>791 </output>
<output>
<ID>OUT_3</ID>781 </output>
<input>
<ID>clear</ID>780 </input>
<input>
<ID>clock</ID>778 </input>
<input>
<ID>count_enable</ID>779 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_REGISTER8</type>
<position>0,13.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>7 </input>
<input>
<ID>IN_4</ID>8 </input>
<input>
<ID>IN_5</ID>9 </input>
<input>
<ID>IN_6</ID>10 </input>
<input>
<ID>IN_7</ID>12 </input>
<input>
<ID>clock</ID>13 </input>
<input>
<ID>load</ID>15 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>781</ID>
<type>AA_TOGGLE</type>
<position>-219.5,-373.5</position>
<output>
<ID>OUT_0</ID>779 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-45.5,-292.5</position>
<gparam>LABEL_TEXT Color Selector Simplified</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>782</ID>
<type>AE_SMALL_INVERTER</type>
<position>-222.5,-378.5</position>
<input>
<ID>IN_0</ID>780 </input>
<output>
<ID>OUT_0</ID>774 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>36.5,29.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>783</ID>
<type>AA_AND2</type>
<position>-217.5,-379.5</position>
<input>
<ID>IN_0</ID>774 </input>
<input>
<ID>IN_1</ID>776 </input>
<output>
<ID>OUT</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_DFF_LOW</type>
<position>53,13</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>55.5,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>59.5,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_OR2</type>
<position>57.5,20</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_DFF_LOW</type>
<position>62,13</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>64.5,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>-26,-27</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>68.5,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_DFF_LOW</type>
<position>-27,-12.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_DFF_LOW</type>
<position>-27,-4</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>-27,4.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_AND2</type>
<position>-195,-354.5</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>795 </input>
<output>
<ID>OUT</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>-27,12.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>795</ID>
<type>AA_TOGGLE</type>
<position>-260,-365</position>
<output>
<ID>OUT_0</ID>796 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>-27,20</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_DFF_LOW</type>
<position>-27,27.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>-27,35</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>10 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_DFF_LOW</type>
<position>-27,42.5</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>799</ID>
<type>AA_LABEL</type>
<position>-263.5,-365</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>-1,6.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-1,21.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>801</ID>
<type>AE_SMALL_INVERTER</type>
<position>-254.5,-365</position>
<input>
<ID>IN_0</ID>796 </input>
<output>
<ID>OUT_0</ID>797 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_OR2</type>
<position>66.5,20</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>802</ID>
<type>AE_SMALL_INVERTER</type>
<position>-250.5,-365</position>
<input>
<ID>IN_0</ID>797 </input>
<output>
<ID>OUT_0</ID>798 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_DFF_LOW</type>
<position>71.5,13</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>803</ID>
<type>AE_SMALL_INVERTER</type>
<position>-235,-365</position>
<input>
<ID>IN_0</ID>798 </input>
<output>
<ID>OUT_0</ID>799 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>74,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>804</ID>
<type>AA_AND2</type>
<position>-227.5,-358.5</position>
<input>
<ID>IN_0</ID>798 </input>
<input>
<ID>IN_1</ID>799 </input>
<output>
<ID>OUT</ID>792 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>-24,56</position>
<gparam>LABEL_TEXT SIPO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>805</ID>
<type>AE_SMALL_INVERTER</type>
<position>-204,-358.5</position>
<input>
<ID>IN_0</ID>792 </input>
<output>
<ID>OUT_0</ID>795 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>78,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_OR2</type>
<position>76,20</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>807</ID>
<type>AE_SMALL_INVERTER</type>
<position>-243.5,-523.5</position>
<input>
<ID>IN_0</ID>801 </input>
<output>
<ID>OUT_0</ID>670 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>80.5,13</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>31 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>808</ID>
<type>AE_SMALL_INVERTER</type>
<position>-243.5,-519.5</position>
<input>
<ID>IN_0</ID>499 </input>
<output>
<ID>OUT_0</ID>801 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>83,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>87,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>810</ID>
<type>AE_SMALL_INVERTER</type>
<position>-37,-536</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>802 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AE_OR2</type>
<position>85,20</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-242.5,-482</position>
<gparam>LABEL_TEXT Change Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>812</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35,-619</position>
<input>
<ID>IN_0</ID>520 </input>
<output>
<ID>OUT_0</ID>803 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>-63.5,-300.5</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>-99,-502.5</position>
<input>
<ID>N_in0</ID>33 </input>
<input>
<ID>N_in1</ID>460 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>168.5,-58.5</position>
<gparam>LABEL_TEXT Notif index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>50.5,-117.5</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>-63,-307</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>-61.5,-304.5</position>
<gparam>LABEL_TEXT Notif Index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>-63,-309</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>-63,-311</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND4</type>
<position>-103,-502.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AI_MUX_8x1</type>
<position>-57.5,-323</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>35 </output>
<input>
<ID>SEL_0</ID>32 </input>
<input>
<ID>SEL_1</ID>29 </input>
<input>
<ID>SEL_2</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>-99,-510.5</position>
<input>
<ID>N_in0</ID>37 </input>
<input>
<ID>N_in1</ID>471 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_MUX_2x1</type>
<position>-31.5,-322.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>53 </output>
<input>
<ID>SEL_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND4</type>
<position>-103,-510.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>91 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>-99,-518.5</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND4</type>
<position>-103,-518.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>92 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>-99,-526.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND4</type>
<position>-103,-526.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>92 </input>
<input>
<ID>IN_3</ID>91 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>-99,-534.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND4</type>
<position>-103,-534.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>89.5,13</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>92,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>96,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR2</type>
<position>94,20</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_DFF_LOW</type>
<position>98.5,13</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>-40.5,-323.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>GA_LED</type>
<position>-99,-542.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND4</type>
<position>-103,-542.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>91 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>101,26</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>105,26</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>103,20</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW</type>
<position>107.5,13</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>clock</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>-99,-550.5</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND4</type>
<position>-103,-550.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>92 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>-99,-558.5</position>
<input>
<ID>N_in0</ID>57 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND4</type>
<position>-103,-558.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>92 </input>
<input>
<ID>IN_3</ID>91 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>24,6.5</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>-66,-325.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>22,20</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>-63,-327</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>-214.5,-550</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>519 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>-20,-322.5</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AE_SMALL_INVERTER</type>
<position>-118,-491.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_SMALL_INVERTER</type>
<position>-114.5,-491.5</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_SMALL_INVERTER</type>
<position>-111,-491.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-40.5,-325</position>
<gparam>LABEL_TEXT Default</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-41,-320.5</position>
<gparam>LABEL_TEXT Custom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>-20,-324.5</position>
<gparam>LABEL_TEXT Light</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>142,-301.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>171.5,-270.5</position>
<gparam>LABEL_TEXT Color Selector</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>138.5,-301.5</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>139.5,-315</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>141,-308.5</position>
<gparam>LABEL_TEXT Notif Index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_TOGGLE</type>
<position>139.5,-313</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>139.5,-311</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>100</ID>
<type>AI_MUX_8x1</type>
<position>144.5,-324</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>73 </output>
<input>
<ID>SEL_0</ID>56 </input>
<input>
<ID>SEL_1</ID>55 </input>
<input>
<ID>SEL_2</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_MUX_2x1</type>
<position>246.5,-328.5</position>
<input>
<ID>IN_0</ID>433 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>421 </output>
<input>
<ID>SEL_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_DFF_LOW</type>
<position>-203,-526</position>
<input>
<ID>IN_0</ID>434 </input>
<output>
<ID>OUT_0</ID>98 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>-200.5,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>-243.5,-535</position>
<input>
<ID>IN_0</ID>670 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>-196.5,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>179.5,-336.5</position>
<gparam>LABEL_TEXT Default</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>58,54.5</position>
<gparam>LABEL_TEXT PISO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>203,-316.5</position>
<gparam>LABEL_TEXT Custom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>300.5,-322</position>
<gparam>LABEL_TEXT Light</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AE_OR2</type>
<position>-198.5,-519</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>437 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_SMALL_INVERTER</type>
<position>-243.5,-539</position>
<input>
<ID>IN_0</ID>530 </input>
<output>
<ID>OUT_0</ID>454 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>-221,-544.5</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>455 </input>
<output>
<ID>OUT</ID>456 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AE_SMALL_INVERTER</type>
<position>-206,-509.5</position>
<input>
<ID>IN_0</ID>570 </input>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_DFF_LOW</type>
<position>-194,-526</position>
<input>
<ID>IN_0</ID>437 </input>
<output>
<ID>OUT_0</ID>144 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_SMALL_INVERTER</type>
<position>-229,-552</position>
<input>
<ID>IN_0</ID>454 </input>
<output>
<ID>OUT_0</ID>455 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>-191.5,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>-187.5,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>449 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>-189.5,-519</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>439 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_DFF_LOW</type>
<position>-185,-526</position>
<input>
<ID>IN_0</ID>439 </input>
<output>
<ID>OUT_0</ID>147 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>-182.5,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>-35.5,-73</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>3,-76</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>-21,-55.5</position>
<gparam>LABEL_TEXT 1:8 Demux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND4</type>
<position>-1,-76</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>85 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>3,-84</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND4</type>
<position>-1,-84</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>104 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>127</ID>
<type>GA_LED</type>
<position>3,-92</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND4</type>
<position>-1,-92</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>85 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>3,-100</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND4</type>
<position>-1,-100</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>104 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>3,-108</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND4</type>
<position>-1,-108</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>85 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>133</ID>
<type>GA_LED</type>
<position>3,-116</position>
<input>
<ID>N_in0</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_AND4</type>
<position>-1,-116</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>86 </input>
<input>
<ID>IN_3</ID>104 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>135</ID>
<type>GA_LED</type>
<position>3,-124</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_AND4</type>
<position>-1,-124</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>85 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>3,-132</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND4</type>
<position>-1,-132</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>106 </input>
<input>
<ID>IN_2</ID>105 </input>
<input>
<ID>IN_3</ID>104 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_TOGGLE</type>
<position>-17.5,-63.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16,-68</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>-14,-63.5</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_SMALL_INVERTER</type>
<position>-12.5,-68</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-63.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AE_SMALL_INVERTER</type>
<position>-9,-68</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>-178.5,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>448 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_DFF_LOW</type>
<position>58,-352</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>60.5,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_OR2</type>
<position>-180.5,-519</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>64.5,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_OR2</type>
<position>62.5,-345</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>46,-345.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_DFF_LOW</type>
<position>-175.5,-526</position>
<input>
<ID>IN_0</ID>438 </input>
<output>
<ID>OUT_0</ID>150 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_SMALL_INVERTER</type>
<position>50.5,-335.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_DFF_LOW</type>
<position>67,-352</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>111 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>-173,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>69.5,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>73.5,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_OR2</type>
<position>71.5,-345</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AE_DFF_LOW</type>
<position>76,-352</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>114 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND2</type>
<position>78.5,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>82.5,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>140 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_OR2</type>
<position>80.5,-345</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_DFF_LOW</type>
<position>85.5,-352</position>
<input>
<ID>IN_0</ID>130 </input>
<output>
<ID>OUT_0</ID>117 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>88,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_AND2</type>
<position>92,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_OR2</type>
<position>90,-345</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_DFF_LOW</type>
<position>94.5,-352</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>120 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND2</type>
<position>97,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND2</type>
<position>101,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_OR2</type>
<position>99,-345</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BB_CLOCK</type>
<position>139,29.5</position>
<output>
<ID>CLK</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>172</ID>
<type>AE_DFF_LOW</type>
<position>103.5,-352</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>123 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>153,32</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>106,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>110,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_OR2</type>
<position>108,-345</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AE_DFF_LOW</type>
<position>112.5,-352</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>126 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>115,-339</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_REGISTER4</type>
<position>151.5,40</position>
<output>
<ID>OUT_3</ID>179 </output>
<input>
<ID>clear</ID>179 </input>
<input>
<ID>clock</ID>177 </input>
<input>
<ID>count_enable</ID>178 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_TOGGLE</type>
<position>144.5,40</position>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_AND2</type>
<position>119,-339</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AE_OR2</type>
<position>117,-345</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_DFF_LOW</type>
<position>121.5,-352</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>359 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>40,-345</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AE_REGISTER8</type>
<position>45,-329.5</position>
<output>
<ID>OUT_0</ID>127 </output>
<output>
<ID>OUT_1</ID>128 </output>
<output>
<ID>OUT_2</ID>141 </output>
<output>
<ID>OUT_3</ID>140 </output>
<output>
<ID>OUT_4</ID>139 </output>
<output>
<ID>OUT_5</ID>138 </output>
<output>
<ID>OUT_6</ID>137 </output>
<output>
<ID>OUT_7</ID>136 </output>
<input>
<ID>clock</ID>153 </input>
<input>
<ID>count_enable</ID>143 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 20</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_SMALL_INVERTER</type>
<position>141.5,35</position>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>44,-336.5</position>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>146.5,34</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_TOGGLE</type>
<position>45,-321.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>-169,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>447 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_OR2</type>
<position>-171,-519</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>440 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AE_DFF_LOW</type>
<position>-166.5,-526</position>
<input>
<ID>IN_0</ID>440 </input>
<output>
<ID>OUT_0</ID>306 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_AND2</type>
<position>-164,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>306 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_AND2</type>
<position>-160,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>446 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_OR2</type>
<position>-162,-519</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>441 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>0.5,-338</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AE_DFF_LOW</type>
<position>56.5,-292.5</position>
<input>
<ID>IN_0</ID>235 </input>
<output>
<ID>OUT_0</ID>160 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>59,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_TOGGLE</type>
<position>137.5,33</position>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_TOGGLE</type>
<position>5.5,-338</position>
<output>
<ID>OUT_0</ID>352 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>63,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_OR2</type>
<position>61,-285.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_TOGGLE</type>
<position>44.5,-286</position>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_OR2</type>
<position>26.5,-336</position>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>353 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AE_OR2</type>
<position>158.5,35</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>49,-276</position>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_DFF_LOW</type>
<position>65.5,-292.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>163 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-343.5</position>
<input>
<ID>IN_0</ID>352 </input>
<output>
<ID>OUT_0</ID>353 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>AE_SMALL_INVERTER</type>
<position>150.5,27.5</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND2</type>
<position>68,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>146,51</position>
<gparam>LABEL_TEXT 8 clock-tick pulse</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AE_DFF_LOW</type>
<position>277.5,6</position>
<input>
<ID>IN_0</ID>203 </input>
<output>
<ID>OUT_0</ID>184 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>280,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>284,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_OR2</type>
<position>282,13</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>265,13</position>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_SMALL_INVERTER</type>
<position>270,22.5</position>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_DFF_LOW</type>
<position>286.5,6</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>187 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND2</type>
<position>289,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>293,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AE_OR2</type>
<position>291,13</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AE_DFF_LOW</type>
<position>295.5,6</position>
<input>
<ID>IN_0</ID>207 </input>
<output>
<ID>OUT_0</ID>190 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND2</type>
<position>298,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND2</type>
<position>302,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_OR2</type>
<position>300,13</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AE_DFF_LOW</type>
<position>305,6</position>
<input>
<ID>IN_0</ID>206 </input>
<output>
<ID>OUT_0</ID>193 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>307.5,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_AND2</type>
<position>311.5,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>AE_OR2</type>
<position>309.5,13</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_DFF_LOW</type>
<position>314,6</position>
<input>
<ID>IN_0</ID>208 </input>
<output>
<ID>OUT_0</ID>196 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>316.5,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_AND2</type>
<position>320.5,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AE_OR2</type>
<position>318.5,13</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>194 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AE_DFF_LOW</type>
<position>323,6</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>199 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_AND2</type>
<position>325.5,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>329.5,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_OR2</type>
<position>327.5,13</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_DFF_LOW</type>
<position>332,6</position>
<input>
<ID>IN_0</ID>210 </input>
<output>
<ID>OUT_0</ID>202 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>334.5,19</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>338.5,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_OR2</type>
<position>336.5,13</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_DFF_LOW</type>
<position>341,6</position>
<input>
<ID>IN_0</ID>211 </input>
<output>
<ID>OUT_0</ID>221 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>72,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>346 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>259.5,13</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AE_OR2</type>
<position>70,-285.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AE_REGISTER8</type>
<position>264.5,28.5</position>
<output>
<ID>OUT_0</ID>203 </output>
<output>
<ID>OUT_1</ID>204 </output>
<output>
<ID>OUT_2</ID>217 </output>
<output>
<ID>OUT_3</ID>216 </output>
<output>
<ID>OUT_4</ID>215 </output>
<output>
<ID>OUT_5</ID>214 </output>
<output>
<ID>OUT_6</ID>213 </output>
<output>
<ID>OUT_7</ID>212 </output>
<input>
<ID>clock</ID>220 </input>
<input>
<ID>count_enable</ID>218 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 37</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_TOGGLE</type>
<position>263.5,21.5</position>
<output>
<ID>OUT_0</ID>220 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>264.5,36.5</position>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_DFF_LOW</type>
<position>74.5,-292.5</position>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>166 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>250</ID>
<type>AE_REGISTER8</type>
<position>403,16</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>223 </input>
<input>
<ID>IN_2</ID>224 </input>
<input>
<ID>IN_3</ID>225 </input>
<input>
<ID>IN_4</ID>226 </input>
<input>
<ID>IN_5</ID>227 </input>
<input>
<ID>IN_6</ID>228 </input>
<input>
<ID>IN_7</ID>230 </input>
<input>
<ID>clock</ID>252 </input>
<input>
<ID>load</ID>232 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND2</type>
<position>77,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>AE_DFF_LOW</type>
<position>376,-10</position>
<input>
<ID>IN_0</ID>221 </input>
<output>
<ID>OUT_0</ID>222 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_DFF_LOW</type>
<position>376,-1.5</position>
<input>
<ID>IN_0</ID>222 </input>
<output>
<ID>OUT_0</ID>223 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_DFF_LOW</type>
<position>376,7</position>
<input>
<ID>IN_0</ID>223 </input>
<output>
<ID>OUT_0</ID>224 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_DFF_LOW</type>
<position>376,15</position>
<input>
<ID>IN_0</ID>224 </input>
<output>
<ID>OUT_0</ID>225 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_DFF_LOW</type>
<position>376,22.5</position>
<input>
<ID>IN_0</ID>225 </input>
<output>
<ID>OUT_0</ID>226 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>257</ID>
<type>AE_DFF_LOW</type>
<position>376,30</position>
<input>
<ID>IN_0</ID>226 </input>
<output>
<ID>OUT_0</ID>227 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>258</ID>
<type>AE_DFF_LOW</type>
<position>376,37.5</position>
<input>
<ID>IN_0</ID>227 </input>
<output>
<ID>OUT_0</ID>228 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_DFF_LOW</type>
<position>376,45</position>
<input>
<ID>IN_0</ID>228 </input>
<output>
<ID>OUT_0</ID>230 </output>
<input>
<ID>clock</ID>247 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_AND2</type>
<position>81,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>345 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>402,24</position>
<output>
<ID>OUT_0</ID>232 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_OR2</type>
<position>79,-285.5</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_DFF_LOW</type>
<position>84,-292.5</position>
<input>
<ID>IN_0</ID>238 </input>
<output>
<ID>OUT_0</ID>170 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_AND2</type>
<position>86.5,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>90.5,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_OR2</type>
<position>88.5,-285.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_DFF_LOW</type>
<position>93,-292.5</position>
<input>
<ID>IN_0</ID>240 </input>
<output>
<ID>OUT_0</ID>174 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>95.5,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>174 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_AND2</type>
<position>99.5,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>343 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_OR2</type>
<position>97.5,-285.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AE_DFF_LOW</type>
<position>102,-292.5</position>
<input>
<ID>IN_0</ID>241 </input>
<output>
<ID>OUT_0</ID>229 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_AND2</type>
<position>104.5,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_TOGGLE</type>
<position>221,3.5</position>
<output>
<ID>OUT_0</ID>246 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_OR2</type>
<position>242,5</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>248 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>AE_SMALL_INVERTER</type>
<position>234,-2.5</position>
<input>
<ID>IN_0</ID>246 </input>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>108.5,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>342 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>BB_CLOCK</type>
<position>222.5,-0.5</position>
<output>
<ID>CLK</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>236.5,2</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_REGISTER4</type>
<position>235,10</position>
<output>
<ID>OUT_3</ID>251 </output>
<input>
<ID>clear</ID>251 </input>
<input>
<ID>clock</ID>249 </input>
<input>
<ID>count_enable</ID>250 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_TOGGLE</type>
<position>228,10</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>281</ID>
<type>AE_SMALL_INVERTER</type>
<position>225,5</position>
<input>
<ID>IN_0</ID>251 </input>
<output>
<ID>OUT_0</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND2</type>
<position>230,4</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_LABEL</type>
<position>217,3</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>AE_OR2</type>
<position>106.5,-285.5</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>AE_SMALL_INVERTER</type>
<position>402,9</position>
<input>
<ID>IN_0</ID>247 </input>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_DFF_LOW</type>
<position>111,-292.5</position>
<input>
<ID>IN_0</ID>312 </input>
<output>
<ID>OUT_0</ID>234 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>287</ID>
<type>GA_LED</type>
<position>185.5,-74.5</position>
<input>
<ID>N_in0</ID>253 </input>
<input>
<ID>N_in1</ID>318 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND4</type>
<position>181.5,-74.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>261 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>289</ID>
<type>GA_LED</type>
<position>185.5,-82.5</position>
<input>
<ID>N_in0</ID>254 </input>
<input>
<ID>N_in1</ID>330 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>AA_AND4</type>
<position>181.5,-82.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>265 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>291</ID>
<type>GA_LED</type>
<position>185.5,-90.5</position>
<input>
<ID>N_in0</ID>255 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_AND4</type>
<position>181.5,-90.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>261 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>293</ID>
<type>GA_LED</type>
<position>185.5,-98.5</position>
<input>
<ID>N_in0</ID>256 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_AND4</type>
<position>181.5,-98.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>263 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>265 </input>
<output>
<ID>OUT</ID>256 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>295</ID>
<type>GA_LED</type>
<position>185.5,-106.5</position>
<input>
<ID>N_in0</ID>257 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND4</type>
<position>181.5,-106.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>261 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>297</ID>
<type>GA_LED</type>
<position>185.5,-114.5</position>
<input>
<ID>N_in0</ID>258 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND4</type>
<position>181.5,-114.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_2</ID>262 </input>
<input>
<ID>IN_3</ID>265 </input>
<output>
<ID>OUT</ID>258 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>299</ID>
<type>GA_LED</type>
<position>185.5,-122.5</position>
<input>
<ID>N_in0</ID>259 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND4</type>
<position>181.5,-122.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>261 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>301</ID>
<type>GA_LED</type>
<position>185.5,-130.5</position>
<input>
<ID>N_in0</ID>260 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND4</type>
<position>181.5,-130.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_2</ID>266 </input>
<input>
<ID>IN_3</ID>265 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_TOGGLE</type>
<position>165,-62</position>
<output>
<ID>OUT_0</ID>267 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_SMALL_INVERTER</type>
<position>166.5,-66.5</position>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>263 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_TOGGLE</type>
<position>168.5,-62</position>
<output>
<ID>OUT_0</ID>266 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_SMALL_INVERTER</type>
<position>170,-66.5</position>
<input>
<ID>IN_0</ID>266 </input>
<output>
<ID>OUT_0</ID>262 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_TOGGLE</type>
<position>172,-62</position>
<output>
<ID>OUT_0</ID>265 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_SMALL_INVERTER</type>
<position>173.5,-66.5</position>
<input>
<ID>IN_0</ID>265 </input>
<output>
<ID>OUT_0</ID>261 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_DFF_LOW</type>
<position>86,-99</position>
<input>
<ID>IN_0</ID>291 </input>
<output>
<ID>OUT_0</ID>272 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_AND2</type>
<position>88.5,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_TOGGLE</type>
<position>55.5,-118</position>
<output>
<ID>OUT_0</ID>311 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_AND2</type>
<position>92.5,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>292 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AE_OR2</type>
<position>90.5,-92</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_TOGGLE</type>
<position>74,-92.5</position>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>315</ID>
<type>AE_OR2</type>
<position>76.5,-116</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AE_SMALL_INVERTER</type>
<position>78.5,-82.5</position>
<input>
<ID>IN_0</ID>270 </input>
<output>
<ID>OUT_0</ID>271 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>317</ID>
<type>AE_DFF_LOW</type>
<position>95,-99</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>275 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_SMALL_INVERTER</type>
<position>68.5,-123.5</position>
<input>
<ID>IN_0</ID>311 </input>
<output>
<ID>OUT_0</ID>313 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>97.5,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>273 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>101.5,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_AND2</type>
<position>113.5,-279.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_OR2</type>
<position>99.5,-92</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>295 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_DFF_LOW</type>
<position>104,-99</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>278 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_AND2</type>
<position>106.5,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>278 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND2</type>
<position>110.5,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_OR2</type>
<position>108.5,-92</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>276 </input>
<output>
<ID>OUT</ID>294 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AE_DFF_LOW</type>
<position>113.5,-99</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>281 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>116,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>281 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>120,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AE_OR2</type>
<position>118,-92</position>
<input>
<ID>IN_0</ID>280 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>296 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AE_DFF_LOW</type>
<position>122.5,-99</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>284 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_REGISTER8</type>
<position>31,35.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<output>
<ID>OUT_1</ID>51 </output>
<output>
<ID>OUT_2</ID>70 </output>
<output>
<ID>OUT_3</ID>69 </output>
<output>
<ID>OUT_4</ID>68 </output>
<output>
<ID>OUT_5</ID>67 </output>
<output>
<ID>OUT_6</ID>66 </output>
<output>
<ID>OUT_7</ID>65 </output>
<input>
<ID>clock</ID>242 </input>
<input>
<ID>count_enable</ID>71 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 18</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_TOGGLE</type>
<position>30,28.5</position>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>31,43.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_AND2</type>
<position>125,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_AND2</type>
<position>129,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>302 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_OR2</type>
<position>127,-92</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>282 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_DFF_LOW</type>
<position>131.5,-99</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>287 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_AND2</type>
<position>134,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>138,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>301 </input>
<output>
<ID>OUT</ID>286 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AE_OR2</type>
<position>136,-92</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>285 </input>
<output>
<ID>OUT</ID>298 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_DFF_LOW</type>
<position>140.5,-99</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>290 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>143,-86</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_AND2</type>
<position>147,-86</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>300 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AE_OR2</type>
<position>145,-92</position>
<input>
<ID>IN_0</ID>289 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_DFF_LOW</type>
<position>149.5,-99</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>264 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>347</ID>
<type>AA_AND2</type>
<position>117.5,-279.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>338 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_LABEL</type>
<position>68,-92</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AE_OR2</type>
<position>115.5,-285.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_REGISTER8</type>
<position>73,-76.5</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>369 </input>
<input>
<ID>IN_2</ID>367 </input>
<input>
<ID>IN_3</ID>366 </input>
<input>
<ID>IN_4</ID>365 </input>
<input>
<ID>IN_5</ID>364 </input>
<input>
<ID>IN_6</ID>363 </input>
<input>
<ID>IN_7</ID>362 </input>
<output>
<ID>OUT_0</ID>291 </output>
<output>
<ID>OUT_1</ID>292 </output>
<output>
<ID>OUT_2</ID>305 </output>
<output>
<ID>OUT_3</ID>304 </output>
<output>
<ID>OUT_4</ID>303 </output>
<output>
<ID>OUT_5</ID>302 </output>
<output>
<ID>OUT_6</ID>301 </output>
<output>
<ID>OUT_7</ID>300 </output>
<input>
<ID>clock</ID>317 </input>
<input>
<ID>load</ID>370 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 202</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_TOGGLE</type>
<position>72,-83.5</position>
<output>
<ID>OUT_0</ID>317 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>352</ID>
<type>AE_DFF_LOW</type>
<position>-157.5,-526</position>
<input>
<ID>IN_0</ID>441 </input>
<output>
<ID>OUT_0</ID>409 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>353</ID>
<type>BB_CLOCK</type>
<position>57,-121.5</position>
<output>
<ID>CLK</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>71,-119</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_REGISTER4</type>
<position>69.5,-111</position>
<output>
<ID>OUT_3</ID>316 </output>
<input>
<ID>clear</ID>316 </input>
<input>
<ID>clock</ID>314 </input>
<input>
<ID>count_enable</ID>315 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_TOGGLE</type>
<position>62.5,-111</position>
<output>
<ID>OUT_0</ID>315 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>357</ID>
<type>AE_SMALL_INVERTER</type>
<position>59.5,-116</position>
<input>
<ID>IN_0</ID>316 </input>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_AND2</type>
<position>64.5,-117</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>311 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AE_DFF_LOW</type>
<position>120,-292.5</position>
<input>
<ID>IN_0</ID>326 </input>
<output>
<ID>OUT_0</ID>360 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>360</ID>
<type>AE_REGISTER8</type>
<position>228,-98</position>
<input>
<ID>IN_0</ID>319 </input>
<input>
<ID>IN_1</ID>320 </input>
<input>
<ID>IN_2</ID>321 </input>
<input>
<ID>IN_3</ID>322 </input>
<input>
<ID>IN_4</ID>323 </input>
<input>
<ID>IN_5</ID>324 </input>
<input>
<ID>IN_6</ID>325 </input>
<input>
<ID>IN_7</ID>327 </input>
<input>
<ID>clock</ID>328 </input>
<input>
<ID>load</ID>329 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>38.5,-285.5</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>AE_DFF_LOW</type>
<position>201,-124</position>
<input>
<ID>IN_0</ID>318 </input>
<output>
<ID>OUT_0</ID>319 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>363</ID>
<type>AE_DFF_LOW</type>
<position>201,-115.5</position>
<input>
<ID>IN_0</ID>319 </input>
<output>
<ID>OUT_0</ID>320 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>364</ID>
<type>AE_DFF_LOW</type>
<position>201,-107</position>
<input>
<ID>IN_0</ID>320 </input>
<output>
<ID>OUT_0</ID>321 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_DFF_LOW</type>
<position>201,-99</position>
<input>
<ID>IN_0</ID>321 </input>
<output>
<ID>OUT_0</ID>322 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_DFF_LOW</type>
<position>201,-91.5</position>
<input>
<ID>IN_0</ID>322 </input>
<output>
<ID>OUT_0</ID>323 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>367</ID>
<type>AE_DFF_LOW</type>
<position>201,-84</position>
<input>
<ID>IN_0</ID>323 </input>
<output>
<ID>OUT_0</ID>324 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_DFF_LOW</type>
<position>201,-76.5</position>
<input>
<ID>IN_0</ID>324 </input>
<output>
<ID>OUT_0</ID>325 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>369</ID>
<type>AE_DFF_LOW</type>
<position>201,-69</position>
<input>
<ID>IN_0</ID>325 </input>
<output>
<ID>OUT_0</ID>327 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_TOGGLE</type>
<position>227,-105</position>
<output>
<ID>OUT_0</ID>328 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_TOGGLE</type>
<position>227,-90</position>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>372</ID>
<type>AE_REGISTER8</type>
<position>43.5,-270</position>
<output>
<ID>OUT_0</ID>235 </output>
<output>
<ID>OUT_1</ID>236 </output>
<output>
<ID>OUT_2</ID>346 </output>
<output>
<ID>OUT_3</ID>345 </output>
<output>
<ID>OUT_4</ID>344 </output>
<output>
<ID>OUT_5</ID>343 </output>
<output>
<ID>OUT_6</ID>342 </output>
<output>
<ID>OUT_7</ID>338 </output>
<input>
<ID>clock</ID>357 </input>
<input>
<ID>count_enable</ID>347 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 21</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_TOGGLE</type>
<position>42.5,-277</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>374</ID>
<type>AE_REGISTER8</type>
<position>231.5,-174.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>332 </input>
<input>
<ID>IN_2</ID>333 </input>
<input>
<ID>IN_3</ID>334 </input>
<input>
<ID>IN_4</ID>335 </input>
<input>
<ID>IN_5</ID>336 </input>
<input>
<ID>IN_6</ID>337 </input>
<input>
<ID>IN_7</ID>339 </input>
<input>
<ID>clock</ID>340 </input>
<input>
<ID>load</ID>341 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_TOGGLE</type>
<position>43.5,-262</position>
<output>
<ID>OUT_0</ID>347 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>376</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-200.5</position>
<input>
<ID>IN_0</ID>330 </input>
<output>
<ID>OUT_0</ID>331 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>377</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-192</position>
<input>
<ID>IN_0</ID>331 </input>
<output>
<ID>OUT_0</ID>332 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>378</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-183.5</position>
<input>
<ID>IN_0</ID>332 </input>
<output>
<ID>OUT_0</ID>333 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-175.5</position>
<input>
<ID>IN_0</ID>333 </input>
<output>
<ID>OUT_0</ID>334 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-168</position>
<input>
<ID>IN_0</ID>334 </input>
<output>
<ID>OUT_0</ID>335 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>381</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-160.5</position>
<input>
<ID>IN_0</ID>335 </input>
<output>
<ID>OUT_0</ID>336 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-153</position>
<input>
<ID>IN_0</ID>336 </input>
<output>
<ID>OUT_0</ID>337 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-145.5</position>
<input>
<ID>IN_0</ID>337 </input>
<output>
<ID>OUT_0</ID>339 </output>
<input>
<ID>clock</ID>307 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_TOGGLE</type>
<position>230.5,-181.5</position>
<output>
<ID>OUT_0</ID>340 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_TOGGLE</type>
<position>230.5,-166.5</position>
<output>
<ID>OUT_0</ID>341 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>386</ID>
<type>BB_CLOCK</type>
<position>5.5,-341.5</position>
<output>
<ID>CLK</ID>349 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>387</ID>
<type>AA_AND2</type>
<position>21,-339</position>
<input>
<ID>IN_0</ID>351 </input>
<input>
<ID>IN_1</ID>349 </input>
<output>
<ID>OUT</ID>348 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_REGISTER4</type>
<position>19.5,-331</position>
<output>
<ID>OUT_3</ID>356 </output>
<input>
<ID>clear</ID>356 </input>
<input>
<ID>clock</ID>354 </input>
<input>
<ID>count_enable</ID>355 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>389</ID>
<type>AA_TOGGLE</type>
<position>12.5,-331</position>
<output>
<ID>OUT_0</ID>355 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>390</ID>
<type>AE_SMALL_INVERTER</type>
<position>9.5,-336</position>
<input>
<ID>IN_0</ID>356 </input>
<output>
<ID>OUT_0</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_AND2</type>
<position>14.5,-337</position>
<input>
<ID>IN_0</ID>350 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>AA_AND2</type>
<position>-155,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_TOGGLE</type>
<position>54,-70.5</position>
<output>
<ID>OUT_0</ID>362 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_TOGGLE</type>
<position>54,-72.5</position>
<output>
<ID>OUT_0</ID>363 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_TOGGLE</type>
<position>54,-74.5</position>
<output>
<ID>OUT_0</ID>364 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_TOGGLE</type>
<position>54,-76.5</position>
<output>
<ID>OUT_0</ID>365 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_TOGGLE</type>
<position>54,-78.5</position>
<output>
<ID>OUT_0</ID>366 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>398</ID>
<type>AA_TOGGLE</type>
<position>54,-80.5</position>
<output>
<ID>OUT_0</ID>367 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>399</ID>
<type>AA_TOGGLE</type>
<position>54,-82.5</position>
<output>
<ID>OUT_0</ID>369 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>400</ID>
<type>AA_TOGGLE</type>
<position>54,-84.5</position>
<output>
<ID>OUT_0</ID>368 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>401</ID>
<type>AA_TOGGLE</type>
<position>72,-68.5</position>
<output>
<ID>OUT_0</ID>370 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>402</ID>
<type>AA_LABEL</type>
<position>48,-77.5</position>
<gparam>LABEL_TEXT New Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AA_LABEL</type>
<position>-77,-322</position>
<gparam>LABEL_TEXT Stored Custom Colors</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>AE_DFF_LOW</type>
<position>177,-369</position>
<input>
<ID>IN_0</ID>394 </input>
<output>
<ID>OUT_0</ID>375 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>179.5,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>371 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>183.5,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>395 </input>
<output>
<ID>OUT</ID>372 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AE_OR2</type>
<position>181.5,-362</position>
<input>
<ID>IN_0</ID>372 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_TOGGLE</type>
<position>165,-362.5</position>
<output>
<ID>OUT_0</ID>373 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>409</ID>
<type>AE_SMALL_INVERTER</type>
<position>169.5,-352.5</position>
<input>
<ID>IN_0</ID>373 </input>
<output>
<ID>OUT_0</ID>374 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_DFF_LOW</type>
<position>186,-369</position>
<input>
<ID>IN_0</ID>396 </input>
<output>
<ID>OUT_0</ID>378 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_AND2</type>
<position>188.5,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>378 </input>
<output>
<ID>OUT</ID>376 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_AND2</type>
<position>192.5,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>408 </input>
<output>
<ID>OUT</ID>377 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>413</ID>
<type>AE_OR2</type>
<position>190.5,-362</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>398 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>AE_DFF_LOW</type>
<position>195,-369</position>
<input>
<ID>IN_0</ID>398 </input>
<output>
<ID>OUT_0</ID>381 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>415</ID>
<type>AA_AND2</type>
<position>197.5,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_AND2</type>
<position>201.5,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>407 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>AE_OR2</type>
<position>199.5,-362</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-369</position>
<input>
<ID>IN_0</ID>397 </input>
<output>
<ID>OUT_0</ID>384 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>419</ID>
<type>AA_AND2</type>
<position>207,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AA_AND2</type>
<position>211,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>406 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>AE_OR2</type>
<position>209,-362</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>382 </input>
<output>
<ID>OUT</ID>399 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>422</ID>
<type>AE_DFF_LOW</type>
<position>213.5,-369</position>
<input>
<ID>IN_0</ID>399 </input>
<output>
<ID>OUT_0</ID>387 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_AND2</type>
<position>216,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>387 </input>
<output>
<ID>OUT</ID>385 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>424</ID>
<type>AA_AND2</type>
<position>220,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>AE_OR2</type>
<position>218,-362</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>400 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>AE_DFF_LOW</type>
<position>222.5,-369</position>
<input>
<ID>IN_0</ID>400 </input>
<output>
<ID>OUT_0</ID>390 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_AND2</type>
<position>225,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>390 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>428</ID>
<type>AA_AND2</type>
<position>229,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>389 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>429</ID>
<type>AE_OR2</type>
<position>227,-362</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>401 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AE_DFF_LOW</type>
<position>231.5,-369</position>
<input>
<ID>IN_0</ID>401 </input>
<output>
<ID>OUT_0</ID>393 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>431</ID>
<type>AA_AND2</type>
<position>234,-356</position>
<input>
<ID>IN_0</ID>373 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>391 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_AND2</type>
<position>238,-356</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>403 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_OR2</type>
<position>236,-362</position>
<input>
<ID>IN_0</ID>392 </input>
<input>
<ID>IN_1</ID>391 </input>
<output>
<ID>OUT</ID>402 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>AE_DFF_LOW</type>
<position>240.5,-369</position>
<input>
<ID>IN_0</ID>402 </input>
<output>
<ID>OUT_0</ID>433 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>159,-362</position>
<gparam>LABEL_TEXT Load/Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AE_REGISTER8</type>
<position>164,-346.5</position>
<input>
<ID>IN_0</ID>412 </input>
<input>
<ID>IN_1</ID>413 </input>
<input>
<ID>IN_2</ID>414 </input>
<input>
<ID>IN_3</ID>415 </input>
<input>
<ID>IN_4</ID>416 </input>
<input>
<ID>IN_5</ID>418 </input>
<input>
<ID>IN_6</ID>417 </input>
<input>
<ID>IN_7</ID>419 </input>
<output>
<ID>OUT_0</ID>394 </output>
<output>
<ID>OUT_1</ID>395 </output>
<output>
<ID>OUT_2</ID>408 </output>
<output>
<ID>OUT_3</ID>407 </output>
<output>
<ID>OUT_4</ID>406 </output>
<output>
<ID>OUT_5</ID>405 </output>
<output>
<ID>OUT_6</ID>404 </output>
<output>
<ID>OUT_7</ID>403 </output>
<input>
<ID>clock</ID>410 </input>
<input>
<ID>load</ID>420 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>437</ID>
<type>AA_TOGGLE</type>
<position>163,-353.5</position>
<output>
<ID>OUT_0</ID>410 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_TOGGLE</type>
<position>163,-338.5</position>
<output>
<ID>OUT_0</ID>420 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>439</ID>
<type>AA_AND2</type>
<position>-151,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>445 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_TOGGLE</type>
<position>152,-339</position>
<output>
<ID>OUT_0</ID>419 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>441</ID>
<type>AA_TOGGLE</type>
<position>152,-341</position>
<output>
<ID>OUT_0</ID>417 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_TOGGLE</type>
<position>152,-343</position>
<output>
<ID>OUT_0</ID>418 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>443</ID>
<type>AA_TOGGLE</type>
<position>152,-345</position>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_TOGGLE</type>
<position>152,-347</position>
<output>
<ID>OUT_0</ID>415 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_TOGGLE</type>
<position>152,-349</position>
<output>
<ID>OUT_0</ID>414 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>446</ID>
<type>AA_TOGGLE</type>
<position>152,-351</position>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>447</ID>
<type>AA_TOGGLE</type>
<position>152,-353</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>448</ID>
<type>AE_OR2</type>
<position>-153,-519</position>
<input>
<ID>IN_0</ID>361 </input>
<input>
<ID>IN_1</ID>358 </input>
<output>
<ID>OUT</ID>442 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_REGISTER8</type>
<position>289,-322.5</position>
<input>
<ID>IN_0</ID>422 </input>
<input>
<ID>IN_1</ID>423 </input>
<input>
<ID>IN_2</ID>424 </input>
<input>
<ID>IN_3</ID>425 </input>
<input>
<ID>IN_4</ID>426 </input>
<input>
<ID>IN_5</ID>427 </input>
<input>
<ID>IN_6</ID>428 </input>
<input>
<ID>IN_7</ID>430 </input>
<input>
<ID>clock</ID>435 </input>
<input>
<ID>load</ID>432 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>450</ID>
<type>AE_DFF_LOW</type>
<position>-148.5,-526</position>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>431 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>451</ID>
<type>AE_DFF_LOW</type>
<position>262,-348.5</position>
<input>
<ID>IN_0</ID>421 </input>
<output>
<ID>OUT_0</ID>422 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>452</ID>
<type>AE_DFF_LOW</type>
<position>262,-340</position>
<input>
<ID>IN_0</ID>422 </input>
<output>
<ID>OUT_0</ID>423 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>453</ID>
<type>AE_DFF_LOW</type>
<position>262,-331.5</position>
<input>
<ID>IN_0</ID>423 </input>
<output>
<ID>OUT_0</ID>424 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>454</ID>
<type>AE_DFF_LOW</type>
<position>262,-323.5</position>
<input>
<ID>IN_0</ID>424 </input>
<output>
<ID>OUT_0</ID>425 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>455</ID>
<type>AE_DFF_LOW</type>
<position>262,-316</position>
<input>
<ID>IN_0</ID>425 </input>
<output>
<ID>OUT_0</ID>426 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>456</ID>
<type>AE_DFF_LOW</type>
<position>262,-308.5</position>
<input>
<ID>IN_0</ID>426 </input>
<output>
<ID>OUT_0</ID>427 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>457</ID>
<type>AE_DFF_LOW</type>
<position>262,-301</position>
<input>
<ID>IN_0</ID>427 </input>
<output>
<ID>OUT_0</ID>428 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>458</ID>
<type>AE_DFF_LOW</type>
<position>262,-293.5</position>
<input>
<ID>IN_0</ID>428 </input>
<output>
<ID>OUT_0</ID>430 </output>
<input>
<ID>clock</ID>348 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>459</ID>
<type>AA_AND2</type>
<position>-146,-513</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_TOGGLE</type>
<position>288,-314.5</position>
<output>
<ID>OUT_0</ID>432 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_AND2</type>
<position>-142,-513</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>444 </input>
<output>
<ID>OUT</ID>429 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_OR2</type>
<position>-144,-519</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>411 </input>
<output>
<ID>OUT</ID>443 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_SMALL_INVERTER</type>
<position>288,-329.5</position>
<input>
<ID>IN_0</ID>348 </input>
<output>
<ID>OUT_0</ID>435 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>465</ID>
<type>AE_DFF_LOW</type>
<position>-139.5,-526</position>
<input>
<ID>IN_0</ID>443 </input>
<output>
<ID>OUT_0</ID>90 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_REGISTER8</type>
<position>-216,-503.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>489 </input>
<input>
<ID>IN_2</ID>487 </input>
<input>
<ID>IN_3</ID>486 </input>
<input>
<ID>IN_4</ID>485 </input>
<input>
<ID>IN_5</ID>484 </input>
<input>
<ID>IN_6</ID>483 </input>
<input>
<ID>IN_7</ID>482 </input>
<output>
<ID>OUT_0</ID>434 </output>
<output>
<ID>OUT_1</ID>436 </output>
<output>
<ID>OUT_2</ID>449 </output>
<output>
<ID>OUT_3</ID>448 </output>
<output>
<ID>OUT_4</ID>447 </output>
<output>
<ID>OUT_5</ID>446 </output>
<output>
<ID>OUT_6</ID>445 </output>
<output>
<ID>OUT_7</ID>444 </output>
<input>
<ID>clock</ID>535 </input>
<input>
<ID>load</ID>490 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>469</ID>
<type>BB_CLOCK</type>
<position>-242,-550</position>
<output>
<ID>CLK</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_AND2</type>
<position>-226.5,-547.5</position>
<input>
<ID>IN_0</ID>453 </input>
<input>
<ID>IN_1</ID>451 </input>
<output>
<ID>OUT</ID>519 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_REGISTER4</type>
<position>-228,-539.5</position>
<output>
<ID>OUT_0</ID>491 </output>
<output>
<ID>OUT_3</ID>459 </output>
<input>
<ID>clear</ID>458 </input>
<input>
<ID>clock</ID>456 </input>
<input>
<ID>count_enable</ID>457 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_TOGGLE</type>
<position>-235,-539.5</position>
<output>
<ID>OUT_0</ID>457 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>473</ID>
<type>AE_SMALL_INVERTER</type>
<position>-238,-544.5</position>
<input>
<ID>IN_0</ID>458 </input>
<output>
<ID>OUT_0</ID>452 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>474</ID>
<type>AA_AND2</type>
<position>-233,-545.5</position>
<input>
<ID>IN_0</ID>452 </input>
<input>
<ID>IN_1</ID>454 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AE_REGISTER8</type>
<position>-36,-529</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>462 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>464 </input>
<input>
<ID>IN_4</ID>465 </input>
<input>
<ID>IN_5</ID>466 </input>
<input>
<ID>IN_6</ID>467 </input>
<input>
<ID>IN_7</ID>468 </input>
<output>
<ID>OUT_0</ID>650 </output>
<output>
<ID>OUT_1</ID>651 </output>
<output>
<ID>OUT_2</ID>652 </output>
<output>
<ID>OUT_3</ID>653 </output>
<output>
<ID>OUT_4</ID>654 </output>
<output>
<ID>OUT_5</ID>804 </output>
<output>
<ID>OUT_6</ID>656 </output>
<output>
<ID>OUT_7</ID>657 </output>
<input>
<ID>clock</ID>802 </input>
<input>
<ID>load</ID>470 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>476</ID>
<type>AE_DFF_LOW</type>
<position>-63,-555</position>
<input>
<ID>IN_0</ID>460 </input>
<output>
<ID>OUT_0</ID>461 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>477</ID>
<type>AE_DFF_LOW</type>
<position>-63,-546.5</position>
<input>
<ID>IN_0</ID>461 </input>
<output>
<ID>OUT_0</ID>462 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>478</ID>
<type>AE_DFF_LOW</type>
<position>-63,-538</position>
<input>
<ID>IN_0</ID>462 </input>
<output>
<ID>OUT_0</ID>463 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>479</ID>
<type>AE_DFF_LOW</type>
<position>-63,-530</position>
<input>
<ID>IN_0</ID>463 </input>
<output>
<ID>OUT_0</ID>464 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>480</ID>
<type>AE_DFF_LOW</type>
<position>-63,-522.5</position>
<input>
<ID>IN_0</ID>464 </input>
<output>
<ID>OUT_0</ID>465 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>481</ID>
<type>AE_DFF_LOW</type>
<position>-63,-515</position>
<input>
<ID>IN_0</ID>465 </input>
<output>
<ID>OUT_0</ID>466 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>482</ID>
<type>AE_DFF_LOW</type>
<position>-63,-507.5</position>
<input>
<ID>IN_0</ID>466 </input>
<output>
<ID>OUT_0</ID>467 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>483</ID>
<type>AE_DFF_LOW</type>
<position>-63,-500</position>
<input>
<ID>IN_0</ID>467 </input>
<output>
<ID>OUT_0</ID>468 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>485</ID>
<type>AA_TOGGLE</type>
<position>-37,-521</position>
<output>
<ID>OUT_0</ID>470 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>486</ID>
<type>AE_REGISTER8</type>
<position>-34,-612</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>473 </input>
<input>
<ID>IN_2</ID>474 </input>
<input>
<ID>IN_3</ID>475 </input>
<input>
<ID>IN_4</ID>476 </input>
<input>
<ID>IN_5</ID>477 </input>
<input>
<ID>IN_6</ID>478 </input>
<input>
<ID>IN_7</ID>479 </input>
<output>
<ID>OUT_0</ID>658 </output>
<output>
<ID>OUT_1</ID>659 </output>
<output>
<ID>OUT_2</ID>660 </output>
<output>
<ID>OUT_3</ID>661 </output>
<output>
<ID>OUT_4</ID>662 </output>
<output>
<ID>OUT_5</ID>663 </output>
<output>
<ID>OUT_6</ID>664 </output>
<output>
<ID>OUT_7</ID>649 </output>
<input>
<ID>clock</ID>803 </input>
<input>
<ID>load</ID>481 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 128</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_DFF_LOW</type>
<position>-61,-638</position>
<input>
<ID>IN_0</ID>471 </input>
<output>
<ID>OUT_0</ID>472 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_DFF_LOW</type>
<position>-61,-629.5</position>
<input>
<ID>IN_0</ID>472 </input>
<output>
<ID>OUT_0</ID>473 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>489</ID>
<type>AE_DFF_LOW</type>
<position>-61,-621</position>
<input>
<ID>IN_0</ID>473 </input>
<output>
<ID>OUT_0</ID>474 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>490</ID>
<type>AE_DFF_LOW</type>
<position>-61,-613</position>
<input>
<ID>IN_0</ID>474 </input>
<output>
<ID>OUT_0</ID>475 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_DFF_LOW</type>
<position>-61,-605.5</position>
<input>
<ID>IN_0</ID>475 </input>
<output>
<ID>OUT_0</ID>476 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>492</ID>
<type>AE_DFF_LOW</type>
<position>-61,-598</position>
<input>
<ID>IN_0</ID>476 </input>
<output>
<ID>OUT_0</ID>477 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>493</ID>
<type>AE_DFF_LOW</type>
<position>-61,-590.5</position>
<input>
<ID>IN_0</ID>477 </input>
<output>
<ID>OUT_0</ID>478 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>494</ID>
<type>AE_DFF_LOW</type>
<position>-61,-583</position>
<input>
<ID>IN_0</ID>478 </input>
<output>
<ID>OUT_0</ID>479 </output>
<input>
<ID>clock</ID>520 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_AND2</type>
<position>-224,-524</position>
<input>
<ID>IN_0</ID>498 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>496</ID>
<type>AA_TOGGLE</type>
<position>-35,-604</position>
<output>
<ID>OUT_0</ID>481 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>497</ID>
<type>AA_TOGGLE</type>
<position>-235,-497.5</position>
<output>
<ID>OUT_0</ID>482 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>498</ID>
<type>AA_TOGGLE</type>
<position>-235,-499.5</position>
<output>
<ID>OUT_0</ID>483 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_TOGGLE</type>
<position>-235,-501.5</position>
<output>
<ID>OUT_0</ID>484 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>500</ID>
<type>AA_TOGGLE</type>
<position>-235,-503.5</position>
<output>
<ID>OUT_0</ID>485 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_TOGGLE</type>
<position>-235,-505.5</position>
<output>
<ID>OUT_0</ID>486 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>502</ID>
<type>AA_TOGGLE</type>
<position>-235,-507.5</position>
<output>
<ID>OUT_0</ID>487 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_TOGGLE</type>
<position>-235,-509.5</position>
<output>
<ID>OUT_0</ID>489 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>504</ID>
<type>AA_TOGGLE</type>
<position>-235,-511.5</position>
<output>
<ID>OUT_0</ID>488 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>505</ID>
<type>AA_TOGGLE</type>
<position>-217,-495.5</position>
<output>
<ID>OUT_0</ID>490 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_LABEL</type>
<position>-241,-504.5</position>
<gparam>LABEL_TEXT New Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>507</ID>
<type>AA_AND2</type>
<position>-206.5,-549</position>
<input>
<ID>IN_0</ID>498 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AE_OR2</type>
<position>-235.5,-517.5</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>499 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_AND2</type>
<position>-206.5,-557</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>807 </input>
<output>
<ID>OUT</ID>450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_AND2</type>
<position>-197,-543.5</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AE_SMALL_INVERTER</type>
<position>-180.5,-540</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>514</ID>
<type>AI_MUX_8x1</type>
<position>84,-583.5</position>
<input>
<ID>IN_0</ID>806 </input>
<input>
<ID>IN_1</ID>805 </input>
<output>
<ID>OUT</ID>494 </output>
<input>
<ID>SEL_0</ID>91 </input>
<input>
<ID>SEL_1</ID>92 </input>
<input>
<ID>SEL_2</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_MUX_2x1</type>
<position>208.5,-581</position>
<input>
<ID>IN_0</ID>645 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>635 </output>
<input>
<ID>SEL_0</ID>807 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_LABEL</type>
<position>132,-596.5</position>
<gparam>LABEL_TEXT Default</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>517</ID>
<type>AA_LABEL</type>
<position>160.5,-577</position>
<gparam>LABEL_TEXT Custom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>518</ID>
<type>AA_LABEL</type>
<position>258.5,-572</position>
<gparam>LABEL_TEXT Light</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>519</ID>
<type>AE_DFF_LOW</type>
<position>3,-611.5</position>
<input>
<ID>IN_0</ID>658 </input>
<output>
<ID>OUT_0</ID>500 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>520</ID>
<type>AA_AND2</type>
<position>5.5,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>500 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>521</ID>
<type>AA_AND2</type>
<position>9.5,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>659 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>522</ID>
<type>AE_OR2</type>
<position>7.5,-604.5</position>
<input>
<ID>IN_0</ID>497 </input>
<input>
<ID>IN_1</ID>496 </input>
<output>
<ID>OUT</ID>521 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>523</ID>
<type>AA_AND2</type>
<position>-179.5,-543.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>528 </input>
<output>
<ID>OUT</ID>655 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>524</ID>
<type>AE_SMALL_INVERTER</type>
<position>-186,-543.5</position>
<input>
<ID>IN_0</ID>532 </input>
<output>
<ID>OUT_0</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>525</ID>
<type>AE_DFF_LOW</type>
<position>12,-611.5</position>
<input>
<ID>IN_0</ID>521 </input>
<output>
<ID>OUT_0</ID>503 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>526</ID>
<type>AA_AND2</type>
<position>14.5,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>503 </input>
<output>
<ID>OUT</ID>501 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_AND2</type>
<position>18.5,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>660 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>AE_OR2</type>
<position>16.5,-604.5</position>
<input>
<ID>IN_0</ID>502 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>523 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>529</ID>
<type>AE_DFF_LOW</type>
<position>21,-611.5</position>
<input>
<ID>IN_0</ID>523 </input>
<output>
<ID>OUT_0</ID>506 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_AND2</type>
<position>23.5,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>506 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_AND2</type>
<position>27.5,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>661 </input>
<output>
<ID>OUT</ID>505 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>532</ID>
<type>AE_OR2</type>
<position>25.5,-604.5</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>504 </input>
<output>
<ID>OUT</ID>522 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>533</ID>
<type>AE_DFF_LOW</type>
<position>30.5,-611.5</position>
<input>
<ID>IN_0</ID>522 </input>
<output>
<ID>OUT_0</ID>509 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>534</ID>
<type>AA_AND2</type>
<position>33,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>509 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_AND2</type>
<position>37,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>662 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>536</ID>
<type>AE_OR2</type>
<position>35,-604.5</position>
<input>
<ID>IN_0</ID>508 </input>
<input>
<ID>IN_1</ID>507 </input>
<output>
<ID>OUT</ID>524 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AE_DFF_LOW</type>
<position>39.5,-611.5</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>512 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>538</ID>
<type>AA_AND2</type>
<position>42,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>AA_AND2</type>
<position>46,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>663 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>540</ID>
<type>AE_OR2</type>
<position>44,-604.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>525 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>541</ID>
<type>AE_DFF_LOW</type>
<position>48.5,-611.5</position>
<input>
<ID>IN_0</ID>525 </input>
<output>
<ID>OUT_0</ID>515 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>542</ID>
<type>AA_AND2</type>
<position>51,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>543</ID>
<type>AA_AND2</type>
<position>55,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>514 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>544</ID>
<type>AE_OR2</type>
<position>53,-604.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>513 </input>
<output>
<ID>OUT</ID>526 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>545</ID>
<type>AE_DFF_LOW</type>
<position>57.5,-611.5</position>
<input>
<ID>IN_0</ID>526 </input>
<output>
<ID>OUT_0</ID>518 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>546</ID>
<type>AA_AND2</type>
<position>60,-598.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>516 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>547</ID>
<type>AA_AND2</type>
<position>64,-598.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>517 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>548</ID>
<type>AE_OR2</type>
<position>62,-604.5</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>516 </input>
<output>
<ID>OUT</ID>527 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>549</ID>
<type>AE_DFF_LOW</type>
<position>66.5,-611.5</position>
<input>
<ID>IN_0</ID>527 </input>
<output>
<ID>OUT_0</ID>805 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>550</ID>
<type>BB_CLOCK</type>
<position>-220,-512.5</position>
<output>
<ID>CLK</ID>535 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>552</ID>
<type>AA_AND2</type>
<position>-213,-515.5</position>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>570 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>554</ID>
<type>AE_DFF_LOW</type>
<position>1.5,-552</position>
<input>
<ID>IN_0</ID>650 </input>
<output>
<ID>OUT_0</ID>540 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>555</ID>
<type>AA_AND2</type>
<position>4,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>540 </input>
<output>
<ID>OUT</ID>536 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>556</ID>
<type>AA_AND2</type>
<position>90,-626.5</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>575 </input>
<output>
<ID>OUT</ID>572 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>AA_AND2</type>
<position>8,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>651 </input>
<output>
<ID>OUT</ID>537 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>558</ID>
<type>AE_OR2</type>
<position>6,-545</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>536 </input>
<output>
<ID>OUT</ID>561 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>559</ID>
<type>AE_SMALL_INVERTER</type>
<position>79.5,-614.5</position>
<input>
<ID>IN_0</ID>584 </input>
<output>
<ID>OUT_0</ID>582 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>560</ID>
<type>AE_SMALL_INVERTER</type>
<position>79.5,-610.5</position>
<input>
<ID>IN_0</ID>648 </input>
<output>
<ID>OUT_0</ID>584 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>105,-642</position>
<input>
<ID>IN_0</ID>579 </input>
<input>
<ID>IN_1</ID>579 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>AE_DFF_LOW</type>
<position>10.5,-552</position>
<input>
<ID>IN_0</ID>561 </input>
<output>
<ID>OUT_0</ID>543 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>563</ID>
<type>AE_SMALL_INVERTER</type>
<position>75,-629.5</position>
<input>
<ID>IN_0</ID>582 </input>
<output>
<ID>OUT_0</ID>580 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>564</ID>
<type>AA_AND2</type>
<position>13,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>543 </input>
<output>
<ID>OUT</ID>541 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_AND2</type>
<position>17,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>652 </input>
<output>
<ID>OUT</ID>542 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>566</ID>
<type>AE_OR2</type>
<position>15,-545</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>541 </input>
<output>
<ID>OUT</ID>563 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>567</ID>
<type>AE_DFF_LOW</type>
<position>19.5,-552</position>
<input>
<ID>IN_0</ID>563 </input>
<output>
<ID>OUT_0</ID>546 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND2</type>
<position>22,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>546 </input>
<output>
<ID>OUT</ID>544 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>569</ID>
<type>AA_AND2</type>
<position>26,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>653 </input>
<output>
<ID>OUT</ID>545 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>570</ID>
<type>AE_OR2</type>
<position>24,-545</position>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>544 </input>
<output>
<ID>OUT</ID>562 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>AE_DFF_LOW</type>
<position>29,-552</position>
<input>
<ID>IN_0</ID>562 </input>
<output>
<ID>OUT_0</ID>549 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_AND2</type>
<position>31.5,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>549 </input>
<output>
<ID>OUT</ID>547 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>573</ID>
<type>AA_AND2</type>
<position>35.5,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>654 </input>
<output>
<ID>OUT</ID>548 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>AE_OR2</type>
<position>33.5,-545</position>
<input>
<ID>IN_0</ID>548 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>564 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>575</ID>
<type>AE_DFF_LOW</type>
<position>38,-552</position>
<input>
<ID>IN_0</ID>564 </input>
<output>
<ID>OUT_0</ID>552 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>576</ID>
<type>AA_AND2</type>
<position>40.5,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>552 </input>
<output>
<ID>OUT</ID>550 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>577</ID>
<type>AA_AND2</type>
<position>44.5,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>804 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>AE_OR2</type>
<position>42.5,-545</position>
<input>
<ID>IN_0</ID>551 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>565 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>579</ID>
<type>AE_DFF_LOW</type>
<position>47,-552</position>
<input>
<ID>IN_0</ID>565 </input>
<output>
<ID>OUT_0</ID>555 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>580</ID>
<type>AA_AND2</type>
<position>49.5,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>555 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>581</ID>
<type>AA_AND2</type>
<position>53.5,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>656 </input>
<output>
<ID>OUT</ID>554 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>582</ID>
<type>AE_OR2</type>
<position>51.5,-545</position>
<input>
<ID>IN_0</ID>554 </input>
<input>
<ID>IN_1</ID>553 </input>
<output>
<ID>OUT</ID>566 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>583</ID>
<type>AE_DFF_LOW</type>
<position>56,-552</position>
<input>
<ID>IN_0</ID>566 </input>
<output>
<ID>OUT_0</ID>558 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_AND2</type>
<position>58.5,-539</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>558 </input>
<output>
<ID>OUT</ID>556 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_AND2</type>
<position>62.5,-539</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>657 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>586</ID>
<type>AE_OR2</type>
<position>60.5,-545</position>
<input>
<ID>IN_0</ID>557 </input>
<input>
<ID>IN_1</ID>556 </input>
<output>
<ID>OUT</ID>567 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>587</ID>
<type>AE_DFF_LOW</type>
<position>65,-552</position>
<input>
<ID>IN_0</ID>567 </input>
<output>
<ID>OUT_0</ID>806 </output>
<input>
<ID>clock</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>588</ID>
<type>AE_SMALL_INVERTER</type>
<position>75,-633.5</position>
<input>
<ID>IN_0</ID>580 </input>
<output>
<ID>OUT_0</ID>560 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_OR2</type>
<position>97.5,-639</position>
<input>
<ID>IN_0</ID>579 </input>
<input>
<ID>IN_1</ID>568 </input>
<output>
<ID>OUT</ID>569 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>590</ID>
<type>AE_SMALL_INVERTER</type>
<position>89.5,-646.5</position>
<input>
<ID>IN_0</ID>560 </input>
<output>
<ID>OUT_0</ID>568 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>591</ID>
<type>BB_CLOCK</type>
<position>76.5,-644.5</position>
<output>
<ID>CLK</ID>538 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>592</ID>
<type>AA_AND2</type>
<position>92,-642</position>
<input>
<ID>IN_0</ID>559 </input>
<input>
<ID>IN_1</ID>538 </input>
<output>
<ID>OUT</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>593</ID>
<type>AA_REGISTER4</type>
<position>90.5,-634</position>
<output>
<ID>OUT_0</ID>575 </output>
<output>
<ID>OUT_3</ID>573 </output>
<input>
<ID>clear</ID>572 </input>
<input>
<ID>clock</ID>569 </input>
<input>
<ID>count_enable</ID>571 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>594</ID>
<type>AA_TOGGLE</type>
<position>83.5,-634</position>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>595</ID>
<type>AE_SMALL_INVERTER</type>
<position>80.5,-639</position>
<input>
<ID>IN_0</ID>572 </input>
<output>
<ID>OUT_0</ID>539 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_AND2</type>
<position>85.5,-640</position>
<input>
<ID>IN_0</ID>539 </input>
<input>
<ID>IN_1</ID>560 </input>
<output>
<ID>OUT</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AE_DFF_LOW</type>
<position>116.5,-628.5</position>
<input>
<ID>IN_0</ID>610 </input>
<output>
<ID>OUT_0</ID>591 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_AND2</type>
<position>119,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>591 </input>
<output>
<ID>OUT</ID>587 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_AND2</type>
<position>123,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>666 </input>
<output>
<ID>OUT</ID>588 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AE_OR2</type>
<position>121,-621.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>587 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_AND2</type>
<position>104.5,-618.5</position>
<input>
<ID>IN_0</ID>581 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>589 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>604</ID>
<type>AE_DFF_LOW</type>
<position>125.5,-628.5</position>
<input>
<ID>IN_0</ID>612 </input>
<output>
<ID>OUT_0</ID>594 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>605</ID>
<type>AA_AND2</type>
<position>128,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>594 </input>
<output>
<ID>OUT</ID>592 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>606</ID>
<type>AA_AND2</type>
<position>132,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>624 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>607</ID>
<type>AE_OR2</type>
<position>130,-621.5</position>
<input>
<ID>IN_0</ID>593 </input>
<input>
<ID>IN_1</ID>592 </input>
<output>
<ID>OUT</ID>614 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>608</ID>
<type>AE_DFF_LOW</type>
<position>134.5,-628.5</position>
<input>
<ID>IN_0</ID>614 </input>
<output>
<ID>OUT_0</ID>597 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_AND2</type>
<position>137,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>597 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_AND2</type>
<position>141,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>623 </input>
<output>
<ID>OUT</ID>596 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>AE_OR2</type>
<position>139,-621.5</position>
<input>
<ID>IN_0</ID>596 </input>
<input>
<ID>IN_1</ID>595 </input>
<output>
<ID>OUT</ID>613 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>612</ID>
<type>AE_DFF_LOW</type>
<position>144,-628.5</position>
<input>
<ID>IN_0</ID>613 </input>
<output>
<ID>OUT_0</ID>600 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_AND2</type>
<position>146.5,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>600 </input>
<output>
<ID>OUT</ID>598 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>614</ID>
<type>AA_AND2</type>
<position>150.5,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>622 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AE_OR2</type>
<position>148.5,-621.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>598 </input>
<output>
<ID>OUT</ID>615 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>616</ID>
<type>AE_DFF_LOW</type>
<position>153,-628.5</position>
<input>
<ID>IN_0</ID>615 </input>
<output>
<ID>OUT_0</ID>603 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_AND2</type>
<position>155.5,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>603 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_AND2</type>
<position>159.5,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>621 </input>
<output>
<ID>OUT</ID>602 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>619</ID>
<type>AE_OR2</type>
<position>157.5,-621.5</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>601 </input>
<output>
<ID>OUT</ID>616 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>620</ID>
<type>AE_DFF_LOW</type>
<position>162,-628.5</position>
<input>
<ID>IN_0</ID>616 </input>
<output>
<ID>OUT_0</ID>606 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>621</ID>
<type>AA_AND2</type>
<position>164.5,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>604 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>622</ID>
<type>AA_AND2</type>
<position>168.5,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>620 </input>
<output>
<ID>OUT</ID>605 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>623</ID>
<type>AE_OR2</type>
<position>166.5,-621.5</position>
<input>
<ID>IN_0</ID>605 </input>
<input>
<ID>IN_1</ID>604 </input>
<output>
<ID>OUT</ID>617 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>624</ID>
<type>AE_DFF_LOW</type>
<position>171,-628.5</position>
<input>
<ID>IN_0</ID>617 </input>
<output>
<ID>OUT_0</ID>609 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>625</ID>
<type>AA_AND2</type>
<position>173.5,-615.5</position>
<input>
<ID>IN_0</ID>589 </input>
<input>
<ID>IN_1</ID>609 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>626</ID>
<type>AA_AND2</type>
<position>177.5,-615.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>619 </input>
<output>
<ID>OUT</ID>608 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_OR2</type>
<position>175.5,-621.5</position>
<input>
<ID>IN_0</ID>608 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>618 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_DFF_LOW</type>
<position>180,-628.5</position>
<input>
<ID>IN_0</ID>618 </input>
<output>
<ID>OUT_0</ID>645 </output>
<input>
<ID>clock</ID>586 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>629</ID>
<type>AE_SMALL_INVERTER</type>
<position>80.5,-620.5</position>
<input>
<ID>IN_0</ID>582 </input>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>630</ID>
<type>AE_REGISTER8</type>
<position>103.5,-606</position>
<input>
<ID>IN_0</ID>626 </input>
<input>
<ID>IN_1</ID>627 </input>
<input>
<ID>IN_2</ID>628 </input>
<input>
<ID>IN_3</ID>629 </input>
<input>
<ID>IN_4</ID>630 </input>
<input>
<ID>IN_5</ID>632 </input>
<input>
<ID>IN_6</ID>631 </input>
<input>
<ID>IN_7</ID>633 </input>
<output>
<ID>OUT_0</ID>610 </output>
<output>
<ID>OUT_1</ID>666 </output>
<output>
<ID>OUT_2</ID>624 </output>
<output>
<ID>OUT_3</ID>623 </output>
<output>
<ID>OUT_4</ID>622 </output>
<output>
<ID>OUT_5</ID>621 </output>
<output>
<ID>OUT_6</ID>620 </output>
<output>
<ID>OUT_7</ID>619 </output>
<input>
<ID>clock</ID>625 </input>
<input>
<ID>load</ID>634 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 135</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>631</ID>
<type>AA_TOGGLE</type>
<position>102.5,-613</position>
<output>
<ID>OUT_0</ID>625 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>632</ID>
<type>AA_TOGGLE</type>
<position>102.5,-598</position>
<output>
<ID>OUT_0</ID>634 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>633</ID>
<type>AA_TOGGLE</type>
<position>91.5,-598.5</position>
<output>
<ID>OUT_0</ID>633 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>634</ID>
<type>AA_TOGGLE</type>
<position>91.5,-600.5</position>
<output>
<ID>OUT_0</ID>631 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>635</ID>
<type>AA_TOGGLE</type>
<position>91.5,-602.5</position>
<output>
<ID>OUT_0</ID>632 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>636</ID>
<type>AA_TOGGLE</type>
<position>91.5,-604.5</position>
<output>
<ID>OUT_0</ID>630 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>637</ID>
<type>AA_TOGGLE</type>
<position>91.5,-606.5</position>
<output>
<ID>OUT_0</ID>629 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>638</ID>
<type>AA_TOGGLE</type>
<position>91.5,-608.5</position>
<output>
<ID>OUT_0</ID>628 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>639</ID>
<type>AA_TOGGLE</type>
<position>91.5,-610.5</position>
<output>
<ID>OUT_0</ID>627 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>640</ID>
<type>AA_TOGGLE</type>
<position>91.5,-612.5</position>
<output>
<ID>OUT_0</ID>626 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_REGISTER8</type>
<position>251,-573.5</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>638 </input>
<input>
<ID>IN_3</ID>639 </input>
<input>
<ID>IN_4</ID>640 </input>
<input>
<ID>IN_5</ID>641 </input>
<input>
<ID>IN_6</ID>642 </input>
<input>
<ID>IN_7</ID>643 </input>
<input>
<ID>clock</ID>667 </input>
<input>
<ID>load</ID>644 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 128</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>642</ID>
<type>AE_DFF_LOW</type>
<position>224,-599.5</position>
<input>
<ID>IN_0</ID>635 </input>
<output>
<ID>OUT_0</ID>636 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>643</ID>
<type>AE_DFF_LOW</type>
<position>224,-591</position>
<input>
<ID>IN_0</ID>636 </input>
<output>
<ID>OUT_0</ID>637 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>644</ID>
<type>AE_DFF_LOW</type>
<position>224,-582.5</position>
<input>
<ID>IN_0</ID>637 </input>
<output>
<ID>OUT_0</ID>638 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_DFF_LOW</type>
<position>224,-574.5</position>
<input>
<ID>IN_0</ID>638 </input>
<output>
<ID>OUT_0</ID>639 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_DFF_LOW</type>
<position>224,-567</position>
<input>
<ID>IN_0</ID>639 </input>
<output>
<ID>OUT_0</ID>640 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_DFF_LOW</type>
<position>224,-559.5</position>
<input>
<ID>IN_0</ID>640 </input>
<output>
<ID>OUT_0</ID>641 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>648</ID>
<type>AE_DFF_LOW</type>
<position>224,-552</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>642 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_DFF_LOW</type>
<position>224,-544.5</position>
<input>
<ID>IN_0</ID>642 </input>
<output>
<ID>OUT_0</ID>643 </output>
<input>
<ID>clock</ID>665 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>650</ID>
<type>AA_TOGGLE</type>
<position>250,-565.5</position>
<output>
<ID>OUT_0</ID>644 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>651</ID>
<type>AE_SMALL_INVERTER</type>
<position>250,-580.5</position>
<input>
<ID>IN_0</ID>665 </input>
<output>
<ID>OUT_0</ID>667 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_AND2</type>
<position>85.5,-619.5</position>
<input>
<ID>IN_0</ID>582 </input>
<input>
<ID>IN_1</ID>583 </input>
<output>
<ID>OUT</ID>576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>653</ID>
<type>AE_SMALL_INVERTER</type>
<position>99.5,-619.5</position>
<input>
<ID>IN_0</ID>576 </input>
<output>
<ID>OUT_0</ID>581 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>655</ID>
<type>AE_SMALL_INVERTER</type>
<position>111,-611.5</position>
<input>
<ID>IN_0</ID>581 </input>
<output>
<ID>OUT_0</ID>647 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_TOGGLE</type>
<position>-235.5,-479.5</position>
<output>
<ID>OUT_0</ID>807 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_TOGGLE</type>
<position>-235.5,-485.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_TOGGLE</type>
<position>-235.5,-487.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>661</ID>
<type>AA_TOGGLE</type>
<position>-235.5,-489.5</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>663</ID>
<type>AA_LABEL</type>
<position>-239,-479.5</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>664</ID>
<type>AA_LABEL</type>
<position>-242,-487.5</position>
<gparam>LABEL_TEXT Notif Index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>665</ID>
<type>AE_SMALL_INVERTER</type>
<position>85.5,-608.5</position>
<input>
<ID>IN_0</ID>807 </input>
<output>
<ID>OUT_0</ID>648 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>667</ID>
<type>AE_OR2</type>
<position>218.5,-625</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>586 </input>
<output>
<ID>OUT</ID>665 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>669</ID>
<type>GA_LED</type>
<position>-191,-354.5</position>
<input>
<ID>N_in0</ID>668 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>670</ID>
<type>GA_LED</type>
<position>-191,-358.5</position>
<input>
<ID>N_in0</ID>669 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>671</ID>
<type>GA_LED</type>
<position>-191,-381.5</position>
<input>
<ID>N_in0</ID>671 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>690</ID>
<type>AE_SMALL_INVERTER</type>
<position>-238,-526</position>
<input>
<ID>IN_0</ID>670 </input>
<output>
<ID>OUT_0</ID>687 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_AND2</type>
<position>-233,-525</position>
<input>
<ID>IN_0</ID>670 </input>
<input>
<ID>IN_1</ID>687 </input>
<output>
<ID>OUT</ID>480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>698</ID>
<type>AE_SMALL_INVERTER</type>
<position>-219,-516.5</position>
<input>
<ID>IN_0</ID>492 </input>
<output>
<ID>OUT_0</ID>570 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>740</ID>
<type>AA_AND2</type>
<position>-213,-366</position>
<input>
<ID>IN_0</ID>781 </input>
<input>
<ID>IN_1</ID>791 </input>
<output>
<ID>OUT</ID>780 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>741</ID>
<type>AA_AND2</type>
<position>-195,-381.5</position>
<input>
<ID>IN_0</ID>793 </input>
<input>
<ID>IN_1</ID>793 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>744</ID>
<type>AE_SMALL_INVERTER</type>
<position>-245.5,-370</position>
<input>
<ID>IN_0</ID>798 </input>
<output>
<ID>OUT_0</ID>794 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>747</ID>
<type>AE_SMALL_INVERTER</type>
<position>-245.5,-374</position>
<input>
<ID>IN_0</ID>794 </input>
<output>
<ID>OUT_0</ID>776 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>748</ID>
<type>AE_OR2</type>
<position>-205.5,-378.5</position>
<input>
<ID>IN_0</ID>793 </input>
<input>
<ID>IN_1</ID>777 </input>
<output>
<ID>OUT</ID>778 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>749</ID>
<type>AE_SMALL_INVERTER</type>
<position>-194,-358.5</position>
<input>
<ID>IN_0</ID>795 </input>
<output>
<ID>OUT_0</ID>669 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_SMALL_INVERTER</type>
<position>-213.5,-386</position>
<input>
<ID>IN_0</ID>776 </input>
<output>
<ID>OUT_0</ID>777 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46.5,23,47.5,23</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<connection>
<GID>5</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>49.5,23,50.5,23</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-21.5,-29,-15.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42,-21.5,-29,-21.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-230,-383,-214,-383</points>
<connection>
<GID>778</GID>
<name>CLK</name></connection>
<intersection>-214 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-214,-383,-214,-382.5</points>
<connection>
<GID>779</GID>
<name>IN_1</name></connection>
<intersection>-383 3</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-9.5,-29,-7</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-8.5,-6,-8.5</points>
<intersection>-29 0</intersection>
<intersection>-6 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-6,-8.5,-6,10.5</points>
<intersection>-8.5 1</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-6,10.5,-4,10.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-6 2</intersection></hsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220.5,-378.5,-220.5,-378.5</points>
<connection>
<GID>782</GID>
<name>OUT_0</name></connection>
<connection>
<GID>783</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-1,-29,1.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>1.78814e-006 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-29,1.78814e-006,-7,1.78814e-006</points>
<intersection>-29 0</intersection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,1.78814e-006,-7,11.5</points>
<intersection>1.78814e-006 3</intersection>
<intersection>11.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,11.5,-4,11.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-7 4</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-214,-380.5,-214,-379.5</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<intersection>-379.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-214.5,-379.5,-214,-379.5</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<intersection>-214 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,7.5,-29,9.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>8.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-29,8.5,-8,8.5</points>
<intersection>-29 0</intersection>
<intersection>-8 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-8,8.5,-8,12.5</points>
<intersection>8.5 6</intersection>
<intersection>12.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-8,12.5,-4,12.5</points>
<connection>
<GID>12</GID>
<name>IN_2</name></connection>
<intersection>-8 7</intersection></hsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-245.5,-380.5,-220.5,-380.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>-245.5 14</intersection>
<intersection>-221.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-221.5,-386,-221.5,-380.5</points>
<intersection>-386 10</intersection>
<intersection>-380.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-221.5,-386,-215.5,-386</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-221.5 9</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-245.5,-380.5,-245.5,-376</points>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection>
<intersection>-380.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,15.5,-29,17</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-29,16,-9,16</points>
<intersection>-29 0</intersection>
<intersection>-9 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9,13.5,-9,16</points>
<intersection>13.5 5</intersection>
<intersection>16 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9,13.5,-4,13.5</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<intersection>-9 4</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-204.5,-386,-204.5,-381.5</points>
<connection>
<GID>748</GID>
<name>IN_1</name></connection>
<intersection>-386 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,-386,-204.5,-386</points>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection>
<intersection>-204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,14.5,-8,23.5</points>
<intersection>14.5 5</intersection>
<intersection>23.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-8,14.5,-4,14.5</points>
<connection>
<GID>12</GID>
<name>IN_4</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-29,23.5,-8,23.5</points>
<intersection>-29 8</intersection>
<intersection>-8 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-29,23,-29,24.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>23.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,30.5,-29,32</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-29,31,-7,31</points>
<intersection>-29 0</intersection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,15.5,-7,31</points>
<intersection>15.5 5</intersection>
<intersection>31 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,15.5,-4,15.5</points>
<connection>
<GID>12</GID>
<name>IN_5</name></connection>
<intersection>-7 4</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-208.5,-374.5,-205.5,-374.5</points>
<connection>
<GID>780</GID>
<name>clock</name></connection>
<intersection>-205.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-205.5,-375.5,-205.5,-374.5</points>
<connection>
<GID>748</GID>
<name>OUT</name></connection>
<intersection>-374.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,38,-29,39.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-29,38.5,-6,38.5</points>
<intersection>-29 0</intersection>
<intersection>-6 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-6,16.5,-6,38.5</points>
<intersection>16.5 5</intersection>
<intersection>38.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-6,16.5,-4,16.5</points>
<connection>
<GID>12</GID>
<name>IN_6</name></connection>
<intersection>-6 4</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-217.5,-373.5,-217.5,-373.5</points>
<connection>
<GID>780</GID>
<name>count_enable</name></connection>
<connection>
<GID>781</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-25,-19.5,39.5</points>
<intersection>-25 19</intersection>
<intersection>-15.5 18</intersection>
<intersection>-7 17</intersection>
<intersection>1.5 16</intersection>
<intersection>9.5 15</intersection>
<intersection>17 14</intersection>
<intersection>24.5 13</intersection>
<intersection>32 20</intersection>
<intersection>39.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-26,39.5,-19.5,39.5</points>
<connection>
<GID>30</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-26,24.5,-19.5,24.5</points>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-26,17,-19.5,17</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-26,9.5,-19.5,9.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-26,1.5,-19.5,1.5</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-26,-7,-19.5,-7</points>
<connection>
<GID>24</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-26,-15.5,-19.5,-15.5</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-26,-25,-19.5,-25</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-26,32,-19.5,32</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224.5,-378.5,-224.5,-362.5</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-362.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224.5,-362.5,-208.5,-362.5</points>
<intersection>-224.5 0</intersection>
<intersection>-213 3</intersection>
<intersection>-208.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-208.5,-372.5,-208.5,-362.5</points>
<connection>
<GID>780</GID>
<name>clear</name></connection>
<intersection>-362.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-213,-363,-213,-362.5</points>
<connection>
<GID>740</GID>
<name>OUT</name></connection>
<intersection>-362.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,45.5,-29,48</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,48,-4,48</points>
<intersection>-29 0</intersection>
<intersection>-4 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-4,17.5,-4,48</points>
<connection>
<GID>12</GID>
<name>IN_7</name></connection>
<intersection>48 1</intersection></vsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-214.5,-369.5,-214.5,-369</points>
<connection>
<GID>780</GID>
<name>OUT_3</name></connection>
<intersection>-369 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-214.5,-369,-214,-369</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>-214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,8.5,-1,8.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,31,102,31</points>
<intersection>34.5 3</intersection>
<intersection>47.5 2</intersection>
<intersection>56.5 16</intersection>
<intersection>65.5 17</intersection>
<intersection>75 18</intersection>
<intersection>84 19</intersection>
<intersection>93 20</intersection>
<intersection>102 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>47.5,29,47.5,31</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>34.5,19.5,34.5,31</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>19.5 22</intersection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>102,29,102,31</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>56.5,29,56.5,31</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>65.5,29,65.5,31</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>75,29,75,31</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>84,29,84,31</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>93,29,93,31</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>34,19.5,34.5,19.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>34.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,19.5,-1,19.5</points>
<connection>
<GID>12</GID>
<name>load</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,29.5,106,29.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>51.5 21</intersection>
<intersection>60.5 13</intersection>
<intersection>69.5 14</intersection>
<intersection>79 15</intersection>
<intersection>88 17</intersection>
<intersection>97 18</intersection>
<intersection>106 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>60.5,29,60.5,29.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>69.5,29,69.5,29.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>79,29,79,29.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>88,29,88,29.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>97,29,97,29.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>106,29,106,29.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>51.5,29,51.5,29.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,17.5,44,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,17.5,47,17.5</points>
<intersection>44 0</intersection>
<intersection>47 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,29,45.5,29</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,15,47,17.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>55.5,23,56.5,23</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58.5,23,59.5,23</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,17.5,53,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,17.5,56,17.5</points>
<intersection>53 0</intersection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,29,54.5,29</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,15,56,17.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>64.5,23,65.5,23</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>67.5,23,68.5,23</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-211.5,-369.5,-211.5,-369</points>
<connection>
<GID>780</GID>
<name>OUT_0</name></connection>
<intersection>-369 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-212,-369,-211.5,-369</points>
<connection>
<GID>740</GID>
<name>IN_1</name></connection>
<intersection>-211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,17.5,62,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,17.5,65,17.5</points>
<intersection>62 0</intersection>
<intersection>65 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,29,63.5,29</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,15,65,17.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-224.5,-358.5,-206,-358.5</points>
<connection>
<GID>804</GID>
<name>OUT</name></connection>
<connection>
<GID>805</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>74,23,75,23</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<connection>
<GID>35</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198,-382.5,-198,-380.5</points>
<connection>
<GID>741</GID>
<name>IN_1</name></connection>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>-381.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-208,-381.5,-198,-381.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<connection>
<GID>779</GID>
<name>OUT</name></connection>
<intersection>-198 0</intersection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-245.5,-372,-245.5,-372</points>
<connection>
<GID>744</GID>
<name>OUT_0</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>77,23,78,23</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,17.5,71.5,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,17.5,74.5,17.5</points>
<intersection>71.5 0</intersection>
<intersection>74.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,29,73,29</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74.5,15,74.5,17.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-202,-358.5,-202,-353.5</points>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection>
<intersection>-358.5 7</intersection>
<intersection>-355.5 9</intersection>
<intersection>-353.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-202,-358.5,-196,-358.5</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-202 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-202,-353.5,-198,-353.5</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<intersection>-202 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-202,-355.5,-198,-355.5</points>
<connection>
<GID>794</GID>
<name>IN_1</name></connection>
<intersection>-202 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,23,84,23</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-258,-365,-256.5,-365</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-317.5,-58.5,-311</points>
<connection>
<GID>53</GID>
<name>SEL_2</name></connection>
<intersection>-311 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-311,-58.5,-311</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252.5,-365,-252.5,-365</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<connection>
<GID>802</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-317.5,-57.5,-309</points>
<connection>
<GID>53</GID>
<name>SEL_1</name></connection>
<intersection>-309 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-309,-57.5,-309</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-248.5,-365,-237,-365</points>
<connection>
<GID>802</GID>
<name>OUT_0</name></connection>
<intersection>-245.5 14</intersection>
<intersection>-237 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-237,-365,-237,-357.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<intersection>-365 1</intersection>
<intersection>-357.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-237,-357.5,-230.5,-357.5</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-237 7</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-245.5,-368,-245.5,-365</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-365 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>86,23,87,23</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232.5,-365,-232.5,-359.5</points>
<intersection>-365 1</intersection>
<intersection>-359.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233,-365,-232.5,-365</points>
<connection>
<GID>803</GID>
<name>OUT_0</name></connection>
<intersection>-232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-232.5,-359.5,-230.5,-359.5</points>
<connection>
<GID>804</GID>
<name>IN_1</name></connection>
<intersection>-232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,17.5,80.5,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,17.5,83.5,17.5</points>
<intersection>80.5 0</intersection>
<intersection>83.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,29,82,29</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>80.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83.5,15,83.5,17.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-317.5,-56.5,-307</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>-307 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-307,-56.5,-307</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-243.5,-521.5,-243.5,-521.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<connection>
<GID>808</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-502.5,-100,-502.5</points>
<connection>
<GID>45</GID>
<name>N_in0</name></connection>
<connection>
<GID>52</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-534,-37,-534</points>
<connection>
<GID>810</GID>
<name>OUT_0</name></connection>
<connection>
<GID>475</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-323.5,-33.5,-323.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-617,-35,-617</points>
<connection>
<GID>812</GID>
<name>OUT_0</name></connection>
<connection>
<GID>486</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-536,43.5,-527</points>
<connection>
<GID>577</GID>
<name>IN_1</name></connection>
<intersection>-527 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-527,43.5,-527</points>
<connection>
<GID>475</GID>
<name>OUT_5</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-323,-44,-321.5</points>
<intersection>-323 2</intersection>
<intersection>-321.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,-321.5,-33.5,-321.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54.5,-323,-44,-323</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-609.5,76,-586</points>
<intersection>-609.5 1</intersection>
<intersection>-586 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-609.5,76,-609.5</points>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-586,81,-586</points>
<connection>
<GID>514</GID>
<name>IN_1</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-320,-31.5,-300.5</points>
<connection>
<GID>55</GID>
<name>SEL_0</name></connection>
<intersection>-300.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58,-300.5,-31.5,-300.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-587,74.5,-550</points>
<intersection>-587 2</intersection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-550,74.5,-550</points>
<connection>
<GID>587</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-587,81,-587</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-510.5,-100,-510.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-518.5,-100,-518.5</points>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-233.5,-479.5,208.5,-479.5</points>
<connection>
<GID>657</GID>
<name>OUT_0</name></connection>
<intersection>-229.5 13</intersection>
<intersection>208.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>208.5,-578.5,208.5,-479.5</points>
<connection>
<GID>515</GID>
<name>SEL_0</name></connection>
<intersection>-563.5 23</intersection>
<intersection>-479.5 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-229.5,-518.5,-229.5,-479.5</points>
<intersection>-518.5 14</intersection>
<intersection>-479.5 7</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-232.5,-518.5,-211,-518.5</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-229.5 13</intersection>
<intersection>-211 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-211,-558,-211,-518.5</points>
<intersection>-558 19</intersection>
<intersection>-542.5 22</intersection>
<intersection>-518.5 14</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-211,-558,-209.5,-558</points>
<connection>
<GID>510</GID>
<name>IN_1</name></connection>
<intersection>-211 18</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-211,-542.5,-200,-542.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>-211 18</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>89,-563.5,208.5,-563.5</points>
<intersection>89 24</intersection>
<intersection>208.5 10</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>89,-608.5,89,-563.5</points>
<intersection>-608.5 31</intersection>
<intersection>-563.5 23</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>87.5,-608.5,89,-608.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>89 24</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-526.5,-100,-526.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-100,-534.5,-100,-534.5</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>92,23,93,23</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>95,23,96,23</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,17.5,89.5,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,17.5,92.5,17.5</points>
<intersection>89.5 0</intersection>
<intersection>92.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,29,91,29</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,15,92.5,17.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>101,23,102,23</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<connection>
<GID>71</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>104,23,105,23</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,17.5,98.5,29</points>
<intersection>17.5 1</intersection>
<intersection>29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,17.5,101.5,17.5</points>
<intersection>98.5 0</intersection>
<intersection>101.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,29,100,29</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>98.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101.5,15,101.5,17.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-542.5,-100,-542.5</points>
<connection>
<GID>69</GID>
<name>N_in0</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-550.5,-100,-550.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,-325.5,-60.5,-325.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,15,41,32.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,32.5,41,32.5</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,29,49.5,33.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,33.5,49.5,33.5</points>
<connection>
<GID>332</GID>
<name>OUT_1</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-327,-60.5,-326.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-327 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-327,-60.5,-327</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,-322.5,-21,-322.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-318.5,143.5,-311</points>
<connection>
<GID>100</GID>
<name>SEL_2</name></connection>
<intersection>-311 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-311,143.5,-311</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-318.5,144.5,-313</points>
<connection>
<GID>100</GID>
<name>SEL_1</name></connection>
<intersection>-313 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-313,144.5,-313</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-318.5,145.5,-315</points>
<connection>
<GID>100</GID>
<name>SEL_0</name></connection>
<intersection>-315 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-315,145.5,-315</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100,-558.5,-100,-558.5</points>
<connection>
<GID>77</GID>
<name>N_in0</name></connection>
<connection>
<GID>78</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,15,48.5,17</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,15,50,15</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,15,66.5,17</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,15,68.5,15</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,15,57.5,17</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,15,59,15</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,15,76,17</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,15,77.5,15</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,15,85,17</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,15,86.5,15</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,15,94,17</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,15,95.5,15</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,15,103,17</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,15,104.5,15</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,29,104,39.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,39.5,104,39.5</points>
<connection>
<GID>332</GID>
<name>OUT_7</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,29,95,38.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,38.5,95,38.5</points>
<connection>
<GID>332</GID>
<name>OUT_6</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,29,86,37.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,37.5,86,37.5</points>
<connection>
<GID>332</GID>
<name>OUT_5</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,29,77,36.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,36.5,77,36.5</points>
<connection>
<GID>332</GID>
<name>OUT_4</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,29,67.5,35.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,35.5,67.5,35.5</points>
<connection>
<GID>332</GID>
<name>OUT_3</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,29,58.5,34.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,34.5,58.5,34.5</points>
<connection>
<GID>332</GID>
<name>OUT_2</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,41.5,31,41.5</points>
<connection>
<GID>332</GID>
<name>count_enable</name></connection>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,6.5,104.5,6.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>41 34</intersection>
<intersection>50 35</intersection>
<intersection>59 36</intersection>
<intersection>68.5 37</intersection>
<intersection>77.5 38</intersection>
<intersection>86.5 33</intersection>
<intersection>95.5 32</intersection>
<intersection>104.5 31</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>104.5,6.5,104.5,12</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>95.5,6.5,95.5,12</points>
<connection>
<GID>67</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>86.5,6.5,86.5,12</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>41,6.5,41,12</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>50,6.5,50,12</points>
<connection>
<GID>15</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>59,6.5,59,12</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>68.5,6.5,68.5,12</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>77.5,6.5,77.5,12</points>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<intersection>6.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153,-327.5,244.5,-327.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>153 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>153,-327.5,153,-324</points>
<intersection>-327.5 1</intersection>
<intersection>-324 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>147.5,-324,153,-324</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>153 6</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-326,246.5,-301.5</points>
<connection>
<GID>101</GID>
<name>SEL_0</name></connection>
<intersection>-301.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-301.5,246.5,-301.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>246.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-111,-553.5,-111,-493.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>-553.5 13</intersection>
<intersection>-537.5 10</intersection>
<intersection>-521.5 5</intersection>
<intersection>-505.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-505.5,-106,-505.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-111,-521.5,-106,-521.5</points>
<connection>
<GID>58</GID>
<name>IN_3</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-111,-537.5,-106,-537.5</points>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-111 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-111,-553.5,-106,-553.5</points>
<connection>
<GID>76</GID>
<name>IN_3</name></connection>
<intersection>-111 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114.5,-543.5,-114.5,-493.5</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>-543.5 16</intersection>
<intersection>-535.5 11</intersection>
<intersection>-511.5 3</intersection>
<intersection>-503.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-114.5,-503.5,-106,-503.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-114.5,-511.5,-106,-511.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-114.5,-535.5,-106,-535.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-114.5,-543.5,-106,-543.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-76,2,-76</points>
<connection>
<GID>122</GID>
<name>N_in0</name></connection>
<connection>
<GID>124</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-84,2,-84</points>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<connection>
<GID>126</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-92,2,-92</points>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<connection>
<GID>128</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-100,2,-100</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<connection>
<GID>130</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>2,-108,2,-108</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<connection>
<GID>132</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-116,2,-116</points>
<connection>
<GID>133</GID>
<name>N_in0</name></connection>
<connection>
<GID>134</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-124,2,-124</points>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<connection>
<GID>136</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-132,2,-132</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<connection>
<GID>138</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-127,-9,-70</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>-127 13</intersection>
<intersection>-111 10</intersection>
<intersection>-95 5</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-79,-4,-79</points>
<connection>
<GID>124</GID>
<name>IN_3</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-9,-95,-4,-95</points>
<connection>
<GID>128</GID>
<name>IN_3</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-9,-111,-4,-111</points>
<connection>
<GID>132</GID>
<name>IN_3</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-9,-127,-4,-127</points>
<connection>
<GID>136</GID>
<name>IN_3</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-117,-12.5,-70</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>-117 16</intersection>
<intersection>-109 11</intersection>
<intersection>-85 3</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-77,-4,-77</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12.5,-85,-4,-85</points>
<connection>
<GID>126</GID>
<name>IN_2</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-12.5,-109,-4,-109</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-12.5,-117,-4,-117</points>
<connection>
<GID>134</GID>
<name>IN_2</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-99,-16,-70</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-99 7</intersection>
<intersection>-91 5</intersection>
<intersection>-83 3</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-75,-4,-75</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-83,-4,-83</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-91,-4,-91</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-16,-99,-4,-99</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33.5,-73,-4,-73</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-24.5,-129,-24.5,-73</points>
<intersection>-129 15</intersection>
<intersection>-121 17</intersection>
<intersection>-113 18</intersection>
<intersection>-105 19</intersection>
<intersection>-97 20</intersection>
<intersection>-89 21</intersection>
<intersection>-81 16</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-24.5,-129,-4,-129</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-24.5,-81,-4,-81</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-24.5,-121,-4,-121</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-24.5,-113,-4,-113</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-24.5,-105,-4,-105</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-24.5,-97,-4,-97</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-24.5,-89,-4,-89</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-24.5 13</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-118,-525.5,-118,-493.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>-525.5 7</intersection>
<intersection>-517.5 5</intersection>
<intersection>-509.5 3</intersection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-118,-501.5,-106,-501.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-118,-509.5,-106,-509.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118,-517.5,-106,-517.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-118,-525.5,-106,-525.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-118 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-134,-499.5,-106,-499.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-134 29</intersection>
<intersection>-126.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-126.5,-555.5,-126.5,-499.5</points>
<intersection>-555.5 15</intersection>
<intersection>-547.5 17</intersection>
<intersection>-539.5 18</intersection>
<intersection>-531.5 19</intersection>
<intersection>-523.5 20</intersection>
<intersection>-515.5 21</intersection>
<intersection>-507.5 16</intersection>
<intersection>-499.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-126.5,-555.5,-106,-555.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-126.5,-507.5,-106,-507.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-126.5,-547.5,-106,-547.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-126.5,-539.5,-106,-539.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-126.5,-531.5,-106,-531.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-126.5,-523.5,-106,-523.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-126.5,-515.5,-106,-515.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-126.5 13</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>-134,-524,-134,-499.5</points>
<intersection>-524 30</intersection>
<intersection>-499.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>-136.5,-524,-134,-524</points>
<connection>
<GID>465</GID>
<name>OUT_0</name></connection>
<intersection>-134 29</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>20</ID>
<points>-233.5,-489.5,85,-489.5</points>
<connection>
<GID>661</GID>
<name>OUT_0</name></connection>
<intersection>-112.5 21</intersection>
<intersection>-111 34</intersection>
<intersection>-109 32</intersection>
<intersection>85 31</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-112.5,-545.5,-112.5,-489.5</points>
<intersection>-545.5 27</intersection>
<intersection>-529.5 26</intersection>
<intersection>-513.5 25</intersection>
<intersection>-489.5 20</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-112.5,-513.5,-106,-513.5</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>-112.5 21</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-112.5,-529.5,-106,-529.5</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>-112.5 21</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-112.5,-545.5,-106,-545.5</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>-112.5 21</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>85,-578,85,-489.5</points>
<connection>
<GID>514</GID>
<name>SEL_0</name></connection>
<intersection>-489.5 20</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-109,-561.5,-109,-489.5</points>
<intersection>-561.5 33</intersection>
<intersection>-489.5 20</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-109,-561.5,-106,-561.5</points>
<connection>
<GID>78</GID>
<name>IN_3</name></connection>
<intersection>-109 32</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>-111,-489.5,-111,-489.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-489.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>-233.5,-487.5,84,-487.5</points>
<connection>
<GID>660</GID>
<name>OUT_0</name></connection>
<intersection>-116 24</intersection>
<intersection>-114.5 36</intersection>
<intersection>84 37</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-116,-559.5,-116,-487.5</points>
<intersection>-559.5 39</intersection>
<intersection>-551.5 32</intersection>
<intersection>-527.5 30</intersection>
<intersection>-519.5 28</intersection>
<intersection>-487.5 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-116,-519.5,-106,-519.5</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>-116 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-116,-527.5,-106,-527.5</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>-116 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-116,-551.5,-106,-551.5</points>
<connection>
<GID>76</GID>
<name>IN_2</name></connection>
<intersection>-116 24</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>-114.5,-489.5,-114.5,-487.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-487.5 23</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>84,-578,84,-487.5</points>
<connection>
<GID>514</GID>
<name>SEL_1</name></connection>
<intersection>-487.5 23</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-116,-559.5,-106,-559.5</points>
<connection>
<GID>78</GID>
<name>IN_2</name></connection>
<intersection>-116 24</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>22</ID>
<points>-233.5,-485.5,83,-485.5</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>-119.5 23</intersection>
<intersection>-118 36</intersection>
<intersection>83 37</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-119.5,-557.5,-119.5,-485.5</points>
<intersection>-557.5 39</intersection>
<intersection>-549.5 31</intersection>
<intersection>-541.5 29</intersection>
<intersection>-533.5 27</intersection>
<intersection>-485.5 22</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-119.5,-533.5,-106,-533.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-119.5 23</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-119.5,-541.5,-106,-541.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-119.5 23</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-119.5,-549.5,-106,-549.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-119.5 23</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>-118,-489.5,-118,-485.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-485.5 22</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>83,-578,83,-485.5</points>
<connection>
<GID>514</GID>
<name>SEL_2</name></connection>
<intersection>-485.5 22</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>-119.5,-557.5,-106,-557.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>-119.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-200.5,-516,-199.5,-516</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-197.5,-516,-196.5,-516</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>19</ID>
<points>-131.5,-540,-131.5,-495</points>
<intersection>-540 79</intersection>
<intersection>-495 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-131.5,-495,-6,-495</points>
<intersection>-131.5 19</intersection>
<intersection>-6 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>-6,-595,-6,-495</points>
<intersection>-595 47</intersection>
<intersection>-535 69</intersection>
<intersection>-495 24</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>-6,-595,65,-595</points>
<intersection>-6 36</intersection>
<intersection>10.5 77</intersection>
<intersection>19.5 59</intersection>
<intersection>28.5 60</intersection>
<intersection>38 61</intersection>
<intersection>47 63</intersection>
<intersection>56 64</intersection>
<intersection>65 65</intersection></hsegment>
<vsegment>
<ID>59</ID>
<points>19.5,-595.5,19.5,-595</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<vsegment>
<ID>60</ID>
<points>28.5,-595.5,28.5,-595</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>38,-595.5,38,-595</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>47,-595.5,47,-595</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>56,-595.5,56,-595</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<vsegment>
<ID>65</ID>
<points>65,-595.5,65,-595</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<hsegment>
<ID>69</ID>
<points>-6,-535,63.5,-535</points>
<intersection>-6 36</intersection>
<intersection>9 76</intersection>
<intersection>18 75</intersection>
<intersection>27 74</intersection>
<intersection>36.5 73</intersection>
<intersection>45.5 72</intersection>
<intersection>54.5 71</intersection>
<intersection>63.5 70</intersection></hsegment>
<vsegment>
<ID>70</ID>
<points>63.5,-536,63.5,-535</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>71</ID>
<points>54.5,-536,54.5,-535</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>72</ID>
<points>45.5,-536,45.5,-535</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>36.5,-536,36.5,-535</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>27,-536,27,-535</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>18,-536,18,-535</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>9,-536,9,-535</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>-535 69</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>10.5,-595.5,10.5,-595</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>-595 47</intersection></vsegment>
<hsegment>
<ID>79</ID>
<points>-178.5,-540,-131.5,-540</points>
<connection>
<GID>513</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 19</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-203,-521.5,-203,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-203,-521.5,-200,-521.5</points>
<intersection>-203 0</intersection>
<intersection>-200 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-203,-510,-201.5,-510</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>-203 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-200,-524,-200,-521.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-191.5,-516,-190.5,-516</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<connection>
<GID>116</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-188.5,-516,-187.5,-516</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>60.5,-342,61.5,-342</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<connection>
<GID>147</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>63.5,-342,64.5,-342</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-334,116,-334</points>
<intersection>48.5 3</intersection>
<intersection>61.5 2</intersection>
<intersection>70.5 16</intersection>
<intersection>79.5 17</intersection>
<intersection>89 18</intersection>
<intersection>98 19</intersection>
<intersection>107 20</intersection>
<intersection>116 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>61.5,-336,61.5,-334</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-345.5,48.5,-334</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-345.5 22</intersection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>116,-336,116,-334</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>70.5,-336,70.5,-334</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>79.5,-336,79.5,-334</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>89,-336,89,-334</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>98,-336,98,-334</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>107,-336,107,-334</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-334 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>48,-345.5,48.5,-345.5</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>48.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>20</ID>
<points>-10.5,-66,-9,-66</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-10.5 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>-10.5,-135,-10.5,-65.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>-135 24</intersection>
<intersection>-119 27</intersection>
<intersection>-103 26</intersection>
<intersection>-87 25</intersection>
<intersection>-66 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-10.5,-135,-4,-135</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>-10.5 21</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-10.5,-87,-4,-87</points>
<connection>
<GID>126</GID>
<name>IN_3</name></connection>
<intersection>-10.5 21</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-10.5,-103,-4,-103</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>-10.5 21</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-10.5,-119,-4,-119</points>
<connection>
<GID>134</GID>
<name>IN_3</name></connection>
<intersection>-10.5 21</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>-14,-66,-12.5,-66</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-14 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-14,-133,-14,-65.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-133 27</intersection>
<intersection>-125 32</intersection>
<intersection>-101 30</intersection>
<intersection>-93 28</intersection>
<intersection>-66 23</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-14,-133,-4,-133</points>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<intersection>-14 24</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-14,-93,-4,-93</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>-14 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-14,-101,-4,-101</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>-14 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-14,-125,-4,-125</points>
<connection>
<GID>136</GID>
<name>IN_2</name></connection>
<intersection>-14 24</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>22</ID>
<points>-17.5,-66,-16,-66</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-17.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-17.5,-131,-17.5,-65.5</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<intersection>-131 26</intersection>
<intersection>-123 31</intersection>
<intersection>-115 29</intersection>
<intersection>-107 27</intersection>
<intersection>-66 22</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-17.5,-131,-4,-131</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-17.5 23</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-17.5,-107,-4,-107</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-17.5 23</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-17.5,-115,-4,-115</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>-17.5 23</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-17.5,-123,-4,-123</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>-17.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-335.5,120,-335.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>65.5 21</intersection>
<intersection>74.5 13</intersection>
<intersection>83.5 14</intersection>
<intersection>93 15</intersection>
<intersection>102 17</intersection>
<intersection>111 18</intersection>
<intersection>120 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>74.5,-336,74.5,-335.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>83.5,-336,83.5,-335.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>93,-336,93,-335.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>102,-336,102,-335.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>111,-336,111,-335.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>120,-336,120,-335.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>65.5,-336,65.5,-335.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-335.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-347.5,58,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-347.5,61,-347.5</points>
<intersection>58 0</intersection>
<intersection>61 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58,-336,59.5,-336</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>58 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>61,-350,61,-347.5</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>69.5,-342,70.5,-342</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<connection>
<GID>156</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>72.5,-342,73.5,-342</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-347.5,67,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-347.5,70,-347.5</points>
<intersection>67 0</intersection>
<intersection>70 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67,-336,68.5,-336</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>67 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70,-350,70,-347.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>78.5,-342,79.5,-342</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<connection>
<GID>160</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>81.5,-342,82.5,-342</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-347.5,76,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-347.5,79,-347.5</points>
<intersection>76 0</intersection>
<intersection>79 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-336,77.5,-336</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>76 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>79,-350,79,-347.5</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>88,-342,89,-342</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91,-342,92,-342</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>165</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-347.5,85.5,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-347.5,88.5,-347.5</points>
<intersection>85.5 0</intersection>
<intersection>88.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-336,87,-336</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>85.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88.5,-350,88.5,-347.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>97,-342,98,-342</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100,-342,101,-342</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>169</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-347.5,94.5,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94.5,-347.5,97.5,-347.5</points>
<intersection>94.5 0</intersection>
<intersection>97.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-336,96,-336</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>94.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-350,97.5,-347.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106,-342,107,-342</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109,-342,110,-342</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<connection>
<GID>175</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-347.5,103.5,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-347.5,106.5,-347.5</points>
<intersection>103.5 0</intersection>
<intersection>106.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-336,105,-336</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>103.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>106.5,-350,106.5,-347.5</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>115,-342,116,-342</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<connection>
<GID>178</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118,-342,119,-342</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-347.5,112.5,-336</points>
<intersection>-347.5 1</intersection>
<intersection>-336 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-347.5,115.5,-347.5</points>
<intersection>112.5 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-336,114,-336</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-350,115.5,-347.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-347.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-350,55,-332.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-332.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,-332.5,55,-332.5</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-336,63.5,-331.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-331.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-331.5,63.5,-331.5</points>
<connection>
<GID>185</GID>
<name>OUT_1</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-350,62.5,-348</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-350,64,-350</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-350,80.5,-348</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-350,82.5,-350</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-350,71.5,-348</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-350,73,-350</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-350,90,-348</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-350,91.5,-350</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-350,99,-348</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-350,100.5,-350</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-350,108,-348</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-350,109.5,-350</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-350,117,-348</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>-350 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-350,118.5,-350</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-336,118,-325.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>-325.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-325.5,118,-325.5</points>
<connection>
<GID>185</GID>
<name>OUT_7</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-336,109,-326.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>-326.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-326.5,109,-326.5</points>
<connection>
<GID>185</GID>
<name>OUT_6</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-336,100,-327.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>-327.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-327.5,100,-327.5</points>
<connection>
<GID>185</GID>
<name>OUT_5</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-336,91,-328.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>-328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-328.5,91,-328.5</points>
<connection>
<GID>185</GID>
<name>OUT_4</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-336,81.5,-329.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>-329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-329.5,81.5,-329.5</points>
<connection>
<GID>185</GID>
<name>OUT_3</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-336,72.5,-330.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>-330.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-330.5,72.5,-330.5</points>
<connection>
<GID>185</GID>
<name>OUT_2</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>143,29.5,150,29.5</points>
<connection>
<GID>171</GID>
<name>CLK</name></connection>
<intersection>150 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>150,29.5,150,31</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>29.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-323.5,45,-323.5</points>
<connection>
<GID>185</GID>
<name>count_enable</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-194,-521.5,-194,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-194,-521.5,-191,-521.5</points>
<intersection>-194 0</intersection>
<intersection>-191 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-194,-510,-192.5,-510</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-194 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-191,-524,-191,-521.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-182.5,-516,-181.5,-516</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-179.5,-516,-178.5,-516</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-185,-521.5,-185,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-185,-521.5,-182,-521.5</points>
<intersection>-185 0</intersection>
<intersection>-182 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-185,-510,-183.5,-510</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-185 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-182,-524,-182,-521.5</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-173,-516,-172,-516</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<connection>
<GID>155</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-170,-516,-169,-516</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-175.5,-521.5,-175.5,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-175.5,-521.5,-172.5,-521.5</points>
<intersection>-175.5 0</intersection>
<intersection>-172.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-175.5,-510,-174,-510</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>-175.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-172.5,-524,-172.5,-521.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-164,-516,-163,-516</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>193</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-161,-516,-160,-516</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<connection>
<GID>194</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-334.5,44,-334.5</points>
<connection>
<GID>185</GID>
<name>clock</name></connection>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>59,-282.5,60,-282.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<connection>
<GID>198</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,35,143.5,35</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>62,-282.5,63,-282.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<connection>
<GID>201</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,33,150,34</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>34 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>149.5,34,150,34</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-274.5,114.5,-274.5</points>
<intersection>47 3</intersection>
<intersection>60 2</intersection>
<intersection>69 16</intersection>
<intersection>78 17</intersection>
<intersection>87.5 18</intersection>
<intersection>96.5 19</intersection>
<intersection>105.5 20</intersection>
<intersection>114.5 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>60,-276.5,60,-274.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>47,-286,47,-274.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-286 22</intersection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>114.5,-276.5,114.5,-274.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>69,-276.5,69,-274.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>78,-276.5,78,-274.5</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>87.5,-276.5,87.5,-274.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>96.5,-276.5,96.5,-274.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>105.5,-276.5,105.5,-274.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>-274.5 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>46.5,-286,47,-286</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>47 3</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-276,118.5,-276</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>64 21</intersection>
<intersection>73 13</intersection>
<intersection>82 14</intersection>
<intersection>91.5 15</intersection>
<intersection>100.5 17</intersection>
<intersection>109.5 18</intersection>
<intersection>118.5 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>73,-276.5,73,-276</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>82,-276.5,82,-276</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>91.5,-276.5,91.5,-276</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>100.5,-276.5,100.5,-276</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>109.5,-276.5,109.5,-276</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>118.5,-276.5,118.5,-276</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>64,-276.5,64,-276</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-276 1</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-288,56.5,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-288,59.5,-288</points>
<intersection>56.5 0</intersection>
<intersection>59.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-276.5,58,-276.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-290.5,59.5,-288</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>68,-282.5,69,-282.5</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<connection>
<GID>210</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>71,-282.5,72,-282.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<connection>
<GID>243</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-288,65.5,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-288,68.5,-288</points>
<intersection>65.5 0</intersection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-276.5,67,-276.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68.5,-290.5,68.5,-288</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>77,-282.5,78,-282.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<connection>
<GID>251</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80,-282.5,81,-282.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-288,74.5,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-288,77.5,-288</points>
<intersection>74.5 0</intersection>
<intersection>77.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-276.5,76,-276.5</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77.5,-290.5,77.5,-288</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,33,143.5,33</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>142.5 9</intersection>
<intersection>143.5 11</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>142.5,27.5,142.5,33</points>
<intersection>27.5 10</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>142.5,27.5,148.5,27.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>142.5 9</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>143.5,33,143.5,33</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>33 1</intersection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>86.5,-282.5,87.5,-282.5</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<connection>
<GID>264</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>89.5,-282.5,90.5,-282.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<connection>
<GID>265</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-288,84,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-288,87,-288</points>
<intersection>84 0</intersection>
<intersection>87 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-276.5,85.5,-276.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>84 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87,-290.5,87,-288</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,32,157.5,32</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<connection>
<GID>173</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>95.5,-282.5,96.5,-282.5</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<connection>
<GID>268</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>98.5,-282.5,99.5,-282.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-288,93,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-288,96,-288</points>
<intersection>93 0</intersection>
<intersection>96 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-276.5,94.5,-276.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96,-290.5,96,-288</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,27.5,159.5,32</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,27.5,159.5,27.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>104.5,-282.5,105.5,-282.5</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<connection>
<GID>272</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155.5,39,158.5,39</points>
<connection>
<GID>179</GID>
<name>clock</name></connection>
<intersection>158.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158.5,38,158.5,39</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>39 1</intersection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>146.5,40,146.5,40</points>
<connection>
<GID>179</GID>
<name>count_enable</name></connection>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,35,139.5,46</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,46,155.5,46</points>
<intersection>139.5 0</intersection>
<intersection>149.5 5</intersection>
<intersection>155.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>155.5,41,155.5,46</points>
<connection>
<GID>179</GID>
<name>clear</name></connection>
<intersection>46 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>149.5,44,149.5,46</points>
<connection>
<GID>179</GID>
<name>OUT_3</name></connection>
<intersection>46 1</intersection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>280,16,281,16</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<connection>
<GID>213</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>283,16,284,16</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<connection>
<GID>214</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>268,24,335.5,24</points>
<intersection>268 3</intersection>
<intersection>281 2</intersection>
<intersection>290 16</intersection>
<intersection>299 17</intersection>
<intersection>308.5 18</intersection>
<intersection>317.5 19</intersection>
<intersection>326.5 20</intersection>
<intersection>335.5 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>281,22,281,24</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>268,13,268,24</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>13 29</intersection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>335.5,22,335.5,24</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>290,22,290,24</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>299,22,299,24</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>308.5,22,308.5,24</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>317.5,22,317.5,24</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>326.5,22,326.5,24</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>267,13,268,13</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>268 3</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272,22.5,339.5,22.5</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>285 21</intersection>
<intersection>294 13</intersection>
<intersection>303 14</intersection>
<intersection>312.5 15</intersection>
<intersection>321.5 17</intersection>
<intersection>330.5 18</intersection>
<intersection>339.5 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>294,22,294,22.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>303,22,303,22.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>312.5,22,312.5,22.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>321.5,22,321.5,22.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>330.5,22,330.5,22.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>339.5,22,339.5,22.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>285,22,285,22.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,10.5,277.5,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,10.5,280.5,10.5</points>
<intersection>277.5 0</intersection>
<intersection>280.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277.5,22,279,22</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>277.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>280.5,8,280.5,10.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>289,16,290,16</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<connection>
<GID>219</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>292,16,293,16</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>220</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,10.5,286.5,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,10.5,289.5,10.5</points>
<intersection>286.5 0</intersection>
<intersection>289.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>286.5,22,288,22</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>286.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>289.5,8,289.5,10.5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298,16,299,16</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301,16,302,16</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,10.5,295.5,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,10.5,298.5,10.5</points>
<intersection>295.5 0</intersection>
<intersection>298.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>295.5,22,297,22</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>295.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>298.5,8,298.5,10.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>307.5,16,308.5,16</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<connection>
<GID>227</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>310.5,16,311.5,16</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305,10.5,305,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>305,10.5,308,10.5</points>
<intersection>305 0</intersection>
<intersection>308 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305,22,306.5,22</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>305 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>308,8,308,10.5</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>316.5,16,317.5,16</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<connection>
<GID>231</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>319.5,16,320.5,16</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,10.5,314,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,10.5,317,10.5</points>
<intersection>314 0</intersection>
<intersection>317 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314,22,315.5,22</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>314 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>317,8,317,10.5</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>325.5,16,326.5,16</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<connection>
<GID>235</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>328.5,16,329.5,16</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<connection>
<GID>236</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,10.5,323,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,10.5,326,10.5</points>
<intersection>323 0</intersection>
<intersection>326 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>323,22,324.5,22</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>323 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>326,8,326,10.5</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>334.5,16,335.5,16</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<connection>
<GID>239</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>337.5,16,338.5,16</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,10.5,332,22</points>
<intersection>10.5 1</intersection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,10.5,335,10.5</points>
<intersection>332 0</intersection>
<intersection>335 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>332,22,333.5,22</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>335,8,335,10.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,8,274.5,25.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>268.5,25.5,274.5,25.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283,22,283,26.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,26.5,283,26.5</points>
<connection>
<GID>246</GID>
<name>OUT_1</name></connection>
<intersection>283 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,8,282,10</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,8,283.5,8</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300,8,300,10</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300,8,302,8</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>300 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,8,291,10</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>291,8,292.5,8</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,8,309.5,10</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,8,311,8</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,8,318.5,10</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,8,320,8</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,8,327.5,10</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,8,329,8</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,8,336.5,10</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336.5,8,338,8</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>336.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337.5,22,337.5,32.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,32.5,337.5,32.5</points>
<connection>
<GID>246</GID>
<name>OUT_7</name></connection>
<intersection>337.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328.5,22,328.5,31.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,31.5,328.5,31.5</points>
<connection>
<GID>246</GID>
<name>OUT_6</name></connection>
<intersection>328.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,22,319.5,30.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,30.5,319.5,30.5</points>
<connection>
<GID>246</GID>
<name>OUT_5</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310.5,22,310.5,29.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,29.5,310.5,29.5</points>
<connection>
<GID>246</GID>
<name>OUT_4</name></connection>
<intersection>310.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301,22,301,28.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,28.5,301,28.5</points>
<connection>
<GID>246</GID>
<name>OUT_3</name></connection>
<intersection>301 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,22,292,27.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,27.5,292,27.5</points>
<connection>
<GID>246</GID>
<name>OUT_2</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,34.5,264.5,34.5</points>
<connection>
<GID>246</GID>
<name>count_enable</name></connection>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>107.5,-282.5,108.5,-282.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<connection>
<GID>276</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,23.5,263.5,23.5</points>
<connection>
<GID>246</GID>
<name>clock</name></connection>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,-14,374,-13</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,-14,374,-14</points>
<intersection>347 3</intersection>
<intersection>374 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>347,-14,347,8</points>
<intersection>-14 1</intersection>
<intersection>8 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>344,8,347,8</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>347 3</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,-7,374,-4.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374,-6,397,-6</points>
<intersection>374 0</intersection>
<intersection>397 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>397,-6,397,13</points>
<intersection>-6 1</intersection>
<intersection>13 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>397,13,399,13</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>397 2</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,1.5,374,4</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>2.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>374,2.5,396,2.5</points>
<intersection>374 0</intersection>
<intersection>396 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>396,2.5,396,14</points>
<intersection>2.5 3</intersection>
<intersection>14 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>396,14,399,14</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>396 4</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,10,374,12</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>11 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>374,11,395,11</points>
<intersection>374 0</intersection>
<intersection>395 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>395,11,395,15</points>
<intersection>11 6</intersection>
<intersection>15 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>395,15,399,15</points>
<connection>
<GID>250</GID>
<name>IN_2</name></connection>
<intersection>395 7</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,18,374,19.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>18.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>374,18.5,394,18.5</points>
<intersection>374 0</intersection>
<intersection>394 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>394,16,394,18.5</points>
<intersection>16 5</intersection>
<intersection>18.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>394,16,399,16</points>
<connection>
<GID>250</GID>
<name>IN_3</name></connection>
<intersection>394 4</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,17,395,26</points>
<intersection>17 5</intersection>
<intersection>26 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>395,17,399,17</points>
<connection>
<GID>250</GID>
<name>IN_4</name></connection>
<intersection>395 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>374,26,395,26</points>
<intersection>374 8</intersection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>374,25.5,374,27</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>26 6</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,33,374,34.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>33.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>374,33.5,396,33.5</points>
<intersection>374 0</intersection>
<intersection>396 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>396,18,396,33.5</points>
<intersection>18 5</intersection>
<intersection>33.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>396,18,399,18</points>
<connection>
<GID>250</GID>
<name>IN_5</name></connection>
<intersection>396 4</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,40.5,374,42</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>41 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>374,41,397,41</points>
<intersection>374 0</intersection>
<intersection>397 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>397,19,397,41</points>
<intersection>19 5</intersection>
<intersection>41 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>397,19,399,19</points>
<connection>
<GID>250</GID>
<name>IN_6</name></connection>
<intersection>397 4</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-288,102,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-288,105,-288</points>
<intersection>102 0</intersection>
<intersection>105 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-276.5,103.5,-276.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>102 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>105,-290.5,105,-288</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>374,48,374,50.5</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>374,50.5,399,50.5</points>
<intersection>374 0</intersection>
<intersection>399 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>399,20,399,50.5</points>
<connection>
<GID>250</GID>
<name>IN_7</name></connection>
<intersection>50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>113.5,-282.5,114.5,-282.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<connection>
<GID>321</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402,22,402,22</points>
<connection>
<GID>250</GID>
<name>load</name></connection>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>116.5,-282.5,117.5,-282.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-288,111,-276.5</points>
<intersection>-288 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-288,114,-288</points>
<intersection>111 0</intersection>
<intersection>114 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-276.5,112.5,-276.5</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-290.5,114,-288</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-290.5,53.5,-273</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-273 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-273,53.5,-273</points>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-276.5,62,-272</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>-272 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-272,62,-272</points>
<connection>
<GID>372</GID>
<name>OUT_1</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-290.5,61,-288.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-290.5,62.5,-290.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-290.5,79,-288.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-290.5,81,-290.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-290.5,70,-288.5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-290.5,71.5,-290.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-290.5,88.5,-288.5</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-290.5,90,-290.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-290.5,97.5,-288.5</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-290.5,99,-290.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,30.5,30,30.5</points>
<connection>
<GID>332</GID>
<name>clock</name></connection>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>226.5,-0.5,233.5,-0.5</points>
<connection>
<GID>277</GID>
<name>CLK</name></connection>
<intersection>233.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>233.5,-0.5,233.5,1</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>-0.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,5,227,5</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<connection>
<GID>282</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233.5,3,233.5,4</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>233,4,233.5,4</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,3.5,227,3.5</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>226 9</intersection>
<intersection>227 13</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>226,-2.5,226,3.5</points>
<intersection>-2.5 10</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>226,-2.5,232,-2.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>226 9</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>227,3,227,3.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239.5,2,241,2</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>241 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>241,-0.5,241,2</points>
<intersection>-0.5 4</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>241,-0.5,338,-0.5</points>
<intersection>241 2</intersection>
<intersection>274.5 37</intersection>
<intersection>283.5 38</intersection>
<intersection>292.5 39</intersection>
<intersection>302 40</intersection>
<intersection>311 41</intersection>
<intersection>320 36</intersection>
<intersection>329 35</intersection>
<intersection>338 34</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>338,-17,338,5</points>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<intersection>-17 60</intersection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>329,-0.5,329,5</points>
<connection>
<GID>238</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>320,-0.5,320,5</points>
<connection>
<GID>234</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>274.5,-0.5,274.5,5</points>
<connection>
<GID>212</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>283.5,-0.5,283.5,5</points>
<connection>
<GID>218</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>292.5,-0.5,292.5,5</points>
<connection>
<GID>222</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>302,-0.5,302,5</points>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>41</ID>
<points>311,-0.5,311,5</points>
<connection>
<GID>230</GID>
<name>clock</name></connection>
<intersection>-0.5 4</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>383.5,-17,383.5,42</points>
<intersection>-17 60</intersection>
<intersection>-13 61</intersection>
<intersection>-4.5 66</intersection>
<intersection>4 59</intersection>
<intersection>12 58</intersection>
<intersection>19.5 57</intersection>
<intersection>27 56</intersection>
<intersection>34.5 63</intersection>
<intersection>42 55</intersection></vsegment>
<hsegment>
<ID>55</ID>
<points>377,42,383.5,42</points>
<connection>
<GID>259</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>377,27,383.5,27</points>
<connection>
<GID>257</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>57</ID>
<points>377,19.5,383.5,19.5</points>
<connection>
<GID>256</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>377,12,383.5,12</points>
<connection>
<GID>255</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>59</ID>
<points>377,4,383.5,4</points>
<connection>
<GID>254</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>338,-17,402,-17</points>
<intersection>338 34</intersection>
<intersection>383.5 43</intersection>
<intersection>402 69</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>377,-13,383.5,-13</points>
<connection>
<GID>252</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>377,34.5,383.5,34.5</points>
<connection>
<GID>258</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<hsegment>
<ID>66</ID>
<points>377,-4.5,383.5,-4.5</points>
<connection>
<GID>253</GID>
<name>clock</name></connection>
<intersection>383.5 43</intersection></hsegment>
<vsegment>
<ID>69</ID>
<points>402,-17,402,7</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>-17 60</intersection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-2.5,243,2</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-2.5,243,-2.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>243 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>239,9,242,9</points>
<connection>
<GID>279</GID>
<name>clock</name></connection>
<intersection>242 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>242,8,242,9</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>9 1</intersection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>230,10,230,10</points>
<connection>
<GID>279</GID>
<name>count_enable</name></connection>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,5,223,16</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223,16,239,16</points>
<intersection>223 0</intersection>
<intersection>233 5</intersection>
<intersection>239 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>239,11,239,16</points>
<connection>
<GID>279</GID>
<name>clear</name></connection>
<intersection>16 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>233,14,233,16</points>
<connection>
<GID>279</GID>
<name>OUT_3</name></connection>
<intersection>16 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402,11,402,11</points>
<connection>
<GID>250</GID>
<name>clock</name></connection>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-74.5,184.5,-74.5</points>
<connection>
<GID>287</GID>
<name>N_in0</name></connection>
<connection>
<GID>288</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-82.5,184.5,-82.5</points>
<connection>
<GID>289</GID>
<name>N_in0</name></connection>
<connection>
<GID>290</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-90.5,184.5,-90.5</points>
<connection>
<GID>291</GID>
<name>N_in0</name></connection>
<connection>
<GID>292</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-98.5,184.5,-98.5</points>
<connection>
<GID>293</GID>
<name>N_in0</name></connection>
<connection>
<GID>294</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184.5,-106.5,184.5,-106.5</points>
<connection>
<GID>295</GID>
<name>N_in0</name></connection>
<connection>
<GID>296</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-114.5,184.5,-114.5</points>
<connection>
<GID>297</GID>
<name>N_in0</name></connection>
<connection>
<GID>298</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-122.5,184.5,-122.5</points>
<connection>
<GID>299</GID>
<name>N_in0</name></connection>
<connection>
<GID>300</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-130.5,184.5,-130.5</points>
<connection>
<GID>301</GID>
<name>N_in0</name></connection>
<connection>
<GID>302</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-125.5,173.5,-68.5</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<intersection>-125.5 13</intersection>
<intersection>-109.5 10</intersection>
<intersection>-93.5 5</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,-77.5,178.5,-77.5</points>
<connection>
<GID>288</GID>
<name>IN_3</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>173.5,-93.5,178.5,-93.5</points>
<connection>
<GID>292</GID>
<name>IN_3</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>173.5,-109.5,178.5,-109.5</points>
<connection>
<GID>296</GID>
<name>IN_3</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>173.5,-125.5,178.5,-125.5</points>
<connection>
<GID>300</GID>
<name>IN_3</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-115.5,170,-68.5</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<intersection>-115.5 16</intersection>
<intersection>-107.5 11</intersection>
<intersection>-83.5 3</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-75.5,178.5,-75.5</points>
<connection>
<GID>288</GID>
<name>IN_2</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>170,-83.5,178.5,-83.5</points>
<connection>
<GID>290</GID>
<name>IN_2</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>170,-107.5,178.5,-107.5</points>
<connection>
<GID>296</GID>
<name>IN_2</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>170,-115.5,178.5,-115.5</points>
<connection>
<GID>298</GID>
<name>IN_2</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-97.5,166.5,-68.5</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 7</intersection>
<intersection>-89.5 5</intersection>
<intersection>-81.5 3</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-73.5,178.5,-73.5</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>166.5,-81.5,178.5,-81.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>166.5,-89.5,178.5,-89.5</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>166.5,-97.5,178.5,-97.5</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>150.5,-71.5,178.5,-71.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>150.5 29</intersection>
<intersection>158 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>158,-127.5,158,-71.5</points>
<intersection>-127.5 15</intersection>
<intersection>-119.5 17</intersection>
<intersection>-111.5 18</intersection>
<intersection>-103.5 19</intersection>
<intersection>-95.5 20</intersection>
<intersection>-87.5 21</intersection>
<intersection>-79.5 16</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>158,-127.5,178.5,-127.5</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>158,-79.5,178.5,-79.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>158,-119.5,178.5,-119.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>158,-111.5,178.5,-111.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>158,-103.5,178.5,-103.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>158,-95.5,178.5,-95.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>158,-87.5,178.5,-87.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>158 13</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>150.5,-97,150.5,-71.5</points>
<intersection>-97 30</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>150.5,-97,152.5,-97</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>150.5 29</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>20</ID>
<points>172,-64.5,173.5,-64.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>172 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>172,-133.5,172,-64</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>-133.5 24</intersection>
<intersection>-117.5 27</intersection>
<intersection>-101.5 26</intersection>
<intersection>-85.5 25</intersection>
<intersection>-64.5 20</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>172,-133.5,178.5,-133.5</points>
<connection>
<GID>302</GID>
<name>IN_3</name></connection>
<intersection>172 21</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>172,-85.5,178.5,-85.5</points>
<connection>
<GID>290</GID>
<name>IN_3</name></connection>
<intersection>172 21</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>172,-101.5,178.5,-101.5</points>
<connection>
<GID>294</GID>
<name>IN_3</name></connection>
<intersection>172 21</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>172,-117.5,178.5,-117.5</points>
<connection>
<GID>298</GID>
<name>IN_3</name></connection>
<intersection>172 21</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>168.5,-64.5,170,-64.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>168.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>168.5,-131.5,168.5,-64</points>
<connection>
<GID>305</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 27</intersection>
<intersection>-123.5 32</intersection>
<intersection>-99.5 30</intersection>
<intersection>-91.5 28</intersection>
<intersection>-64.5 23</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>168.5,-131.5,178.5,-131.5</points>
<connection>
<GID>302</GID>
<name>IN_2</name></connection>
<intersection>168.5 24</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>168.5,-91.5,178.5,-91.5</points>
<connection>
<GID>292</GID>
<name>IN_2</name></connection>
<intersection>168.5 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>168.5,-99.5,178.5,-99.5</points>
<connection>
<GID>294</GID>
<name>IN_2</name></connection>
<intersection>168.5 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>168.5,-123.5,178.5,-123.5</points>
<connection>
<GID>300</GID>
<name>IN_2</name></connection>
<intersection>168.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<hsegment>
<ID>22</ID>
<points>165,-64.5,166.5,-64.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>165 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>165,-129.5,165,-64</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<intersection>-129.5 26</intersection>
<intersection>-121.5 31</intersection>
<intersection>-113.5 29</intersection>
<intersection>-105.5 27</intersection>
<intersection>-64.5 22</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>165,-129.5,178.5,-129.5</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>165 23</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>165,-105.5,178.5,-105.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>165 23</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>165,-113.5,178.5,-113.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>165 23</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>165,-121.5,178.5,-121.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>165 23</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>88.5,-89,89.5,-89</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<connection>
<GID>310</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91.5,-89,92.5,-89</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<connection>
<GID>312</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-81,144,-81</points>
<intersection>76.5 3</intersection>
<intersection>89.5 2</intersection>
<intersection>98.5 16</intersection>
<intersection>107.5 17</intersection>
<intersection>117 18</intersection>
<intersection>126 19</intersection>
<intersection>135 20</intersection>
<intersection>144 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>89.5,-83,89.5,-81</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-92.5,76.5,-81</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-92.5 22</intersection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>144,-83,144,-81</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>98.5,-83,98.5,-81</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>107.5,-83,107.5,-81</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>117,-83,117,-81</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>126,-83,126,-81</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>135,-83,135,-81</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>76,-92.5,76.5,-92.5</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>76.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,-82.5,148,-82.5</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>93.5 21</intersection>
<intersection>102.5 13</intersection>
<intersection>111.5 14</intersection>
<intersection>121 15</intersection>
<intersection>130 17</intersection>
<intersection>139 18</intersection>
<intersection>148 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>102.5,-83,102.5,-82.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>111.5,-83,111.5,-82.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>121,-83,121,-82.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>130,-83,130,-82.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>139,-83,139,-82.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>148,-83,148,-82.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>93.5,-83,93.5,-82.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>-82.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-94.5,86,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-94.5,89,-94.5</points>
<intersection>86 0</intersection>
<intersection>89 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-83,87.5,-83</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89,-97,89,-94.5</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>97.5,-89,98.5,-89</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<connection>
<GID>319</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100.5,-89,101.5,-89</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<connection>
<GID>320</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-94.5,95,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-94.5,98,-94.5</points>
<intersection>95 0</intersection>
<intersection>98 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95,-83,96.5,-83</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>98,-97,98,-94.5</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>106.5,-89,107.5,-89</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<connection>
<GID>324</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>109.5,-89,110.5,-89</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>325</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-94.5,104,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-94.5,107,-94.5</points>
<intersection>104 0</intersection>
<intersection>107 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-83,105.5,-83</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107,-97,107,-94.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>116,-89,117,-89</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<connection>
<GID>328</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>119,-89,120,-89</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>329</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-94.5,113.5,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-94.5,116.5,-94.5</points>
<intersection>113.5 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-83,115,-83</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>113.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-97,116.5,-94.5</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>125,-89,126,-89</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<connection>
<GID>335</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>128,-89,129,-89</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-94.5,122.5,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-94.5,125.5,-94.5</points>
<intersection>122.5 0</intersection>
<intersection>125.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-83,124,-83</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>125.5,-97,125.5,-94.5</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>134,-89,135,-89</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<connection>
<GID>339</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>137,-89,138,-89</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-94.5,131.5,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-94.5,134.5,-94.5</points>
<intersection>131.5 0</intersection>
<intersection>134.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-83,133,-83</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>131.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-97,134.5,-94.5</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>143,-89,144,-89</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<connection>
<GID>343</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>146,-89,147,-89</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>344</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-94.5,140.5,-83</points>
<intersection>-94.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-94.5,143.5,-94.5</points>
<intersection>140.5 0</intersection>
<intersection>143.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-83,142,-83</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>140.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>143.5,-97,143.5,-94.5</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-94.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-97,80,-79.5</points>
<intersection>-97 4</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>77,-79.5,80,-79.5</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>80,-97,83,-97</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-83,91.5,-78.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>-78.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-78.5,91.5,-78.5</points>
<connection>
<GID>350</GID>
<name>OUT_1</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-97,90.5,-95</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-97,92,-97</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-97,108.5,-95</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-97,110.5,-97</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-97,99.5,-95</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-97,101,-97</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-97,118,-95</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-97,119.5,-97</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-97,127,-95</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-97,128.5,-97</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-97,136,-95</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-97,137.5,-97</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-97,145,-95</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-97,146.5,-97</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-83,146,-72.5</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-72.5,146,-72.5</points>
<connection>
<GID>350</GID>
<name>OUT_7</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-83,137,-73.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-73.5,137,-73.5</points>
<connection>
<GID>350</GID>
<name>OUT_6</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-83,128,-74.5</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-74.5,128,-74.5</points>
<connection>
<GID>350</GID>
<name>OUT_5</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-83,119,-75.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-75.5,119,-75.5</points>
<connection>
<GID>350</GID>
<name>OUT_4</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-83,109.5,-76.5</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-76.5,109.5,-76.5</points>
<connection>
<GID>350</GID>
<name>OUT_3</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-83,100.5,-77.5</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-77.5,100.5,-77.5</points>
<connection>
<GID>350</GID>
<name>OUT_2</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-166.5,-521.5,-166.5,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-166.5,-521.5,-163.5,-521.5</points>
<intersection>-166.5 0</intersection>
<intersection>-163.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-166.5,-510,-165,-510</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>-166.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-163.5,-524,-163.5,-521.5</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-119,146.5,-119</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>83 116</intersection>
<intersection>92 115</intersection>
<intersection>101 114</intersection>
<intersection>110.5 117</intersection>
<intersection>119.5 118</intersection>
<intersection>128.5 119</intersection>
<intersection>130 39</intersection>
<intersection>137.5 120</intersection>
<intersection>146.5 121</intersection></hsegment>
<vsegment>
<ID>39</ID>
<points>130,-136.5,130,-119</points>
<intersection>-136.5 58</intersection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>215.5,-136.5,215.5,-72</points>
<intersection>-136.5 58</intersection>
<intersection>-118.5 102</intersection>
<intersection>-110 103</intersection>
<intersection>-102 104</intersection>
<intersection>-94.5 105</intersection>
<intersection>-87 106</intersection>
<intersection>-79.5 107</intersection>
<intersection>-72 108</intersection></vsegment>
<hsegment>
<ID>58</ID>
<points>130,-136.5,236,-136.5</points>
<intersection>130 39</intersection>
<intersection>202 61</intersection>
<intersection>209.5 93</intersection>
<intersection>215.5 40</intersection>
<intersection>236 62</intersection></hsegment>
<vsegment>
<ID>61</ID>
<points>202,-136.5,202,-127</points>
<connection>
<GID>362</GID>
<name>clock</name></connection>
<intersection>-136.5 58</intersection></vsegment>
<vsegment>
<ID>62</ID>
<points>236,-209,236,-136.5</points>
<intersection>-209 75</intersection>
<intersection>-136.5 58</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>217.5,-209,217.5,-159</points>
<intersection>-209 75</intersection>
<intersection>-205.5 80</intersection>
<intersection>-197 79</intersection>
<intersection>-189 78</intersection>
<intersection>-181.5 77</intersection>
<intersection>-174 76</intersection>
<intersection>-166.5 83</intersection>
<intersection>-159 85</intersection></vsegment>
<hsegment>
<ID>75</ID>
<points>209.5,-209,236,-209</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection>
<intersection>236 62</intersection></hsegment>
<hsegment>
<ID>76</ID>
<points>209.5,-174,217.5,-174</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>209.5,-181.5,217.5,-181.5</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>78</ID>
<points>209.5,-189,217.5,-189</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>79</ID>
<points>209.5,-197,217.5,-197</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>80</ID>
<points>209.5,-205.5,217.5,-205.5</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>209.5,-166.5,217.5,-166.5</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<hsegment>
<ID>85</ID>
<points>209.5,-159,217.5,-159</points>
<intersection>209.5 93</intersection>
<intersection>217.5 63</intersection></hsegment>
<vsegment>
<ID>93</ID>
<points>209.5,-209,209.5,-136.5</points>
<intersection>-209 75</intersection>
<intersection>-205.5 80</intersection>
<intersection>-203.5 94</intersection>
<intersection>-197 79</intersection>
<intersection>-195 95</intersection>
<intersection>-189 78</intersection>
<intersection>-186.5 96</intersection>
<intersection>-181.5 77</intersection>
<intersection>-178.5 97</intersection>
<intersection>-174 76</intersection>
<intersection>-171 98</intersection>
<intersection>-166.5 83</intersection>
<intersection>-163.5 99</intersection>
<intersection>-159 85</intersection>
<intersection>-156 100</intersection>
<intersection>-148.5 101</intersection>
<intersection>-136.5 58</intersection></vsegment>
<hsegment>
<ID>94</ID>
<points>205.5,-203.5,209.5,-203.5</points>
<connection>
<GID>376</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>205.5,-195,209.5,-195</points>
<connection>
<GID>377</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>205.5,-186.5,209.5,-186.5</points>
<connection>
<GID>378</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>97</ID>
<points>205.5,-178.5,209.5,-178.5</points>
<connection>
<GID>379</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>205.5,-171,209.5,-171</points>
<connection>
<GID>380</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>99</ID>
<points>205.5,-163.5,209.5,-163.5</points>
<connection>
<GID>381</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>100</ID>
<points>205.5,-156,209.5,-156</points>
<connection>
<GID>382</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>101</ID>
<points>205.5,-148.5,209.5,-148.5</points>
<connection>
<GID>383</GID>
<name>clock</name></connection>
<intersection>209.5 93</intersection></hsegment>
<hsegment>
<ID>102</ID>
<points>202,-118.5,215.5,-118.5</points>
<connection>
<GID>363</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>103</ID>
<points>202,-110,215.5,-110</points>
<connection>
<GID>364</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>104</ID>
<points>202,-102,215.5,-102</points>
<connection>
<GID>365</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>105</ID>
<points>202,-94.5,215.5,-94.5</points>
<connection>
<GID>366</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>106</ID>
<points>202,-87,215.5,-87</points>
<connection>
<GID>367</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>107</ID>
<points>202,-79.5,215.5,-79.5</points>
<connection>
<GID>368</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<hsegment>
<ID>108</ID>
<points>202,-72,215.5,-72</points>
<connection>
<GID>369</GID>
<name>clock</name></connection>
<intersection>215.5 40</intersection></hsegment>
<vsegment>
<ID>114</ID>
<points>101,-119,101,-100</points>
<connection>
<GID>323</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>92,-119,92,-100</points>
<connection>
<GID>317</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>83,-119,83,-100</points>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>110.5,-119,110.5,-100</points>
<connection>
<GID>327</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>119.5,-119,119.5,-100</points>
<connection>
<GID>331</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>119</ID>
<points>128.5,-119,128.5,-100</points>
<connection>
<GID>338</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>120</ID>
<points>137.5,-119,137.5,-100</points>
<connection>
<GID>342</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment>
<vsegment>
<ID>121</ID>
<points>146.5,-119,146.5,-100</points>
<connection>
<GID>346</GID>
<name>clock</name></connection>
<intersection>-119 1</intersection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>61,-121.5,68,-121.5</points>
<connection>
<GID>353</GID>
<name>CLK</name></connection>
<intersection>68 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>68,-121.5,68,-120</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<intersection>-121.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-116,61.5,-116</points>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-118,68,-117</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-117 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>67.5,-117,68,-117</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57.5,-118,61.5,-118</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>60.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>60.5,-123.5,60.5,-118</points>
<intersection>-123.5 10</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>60.5,-123.5,66.5,-123.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>60.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-290.5,106.5,-288.5</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-290.5,108,-290.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-123.5,77.5,-119</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-123.5,77.5,-123.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-112,76.5,-112</points>
<connection>
<GID>355</GID>
<name>clock</name></connection>
<intersection>76.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-113,76.5,-112</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>64.5,-111,64.5,-111</points>
<connection>
<GID>355</GID>
<name>count_enable</name></connection>
<connection>
<GID>356</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-116,57.5,-105</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-105,73.5,-105</points>
<intersection>57.5 0</intersection>
<intersection>67.5 5</intersection>
<intersection>73.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>73.5,-110,73.5,-105</points>
<connection>
<GID>355</GID>
<name>clear</name></connection>
<intersection>-105 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>67.5,-107,67.5,-105</points>
<connection>
<GID>355</GID>
<name>OUT_3</name></connection>
<intersection>-105 1</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-81.5,72,-81.5</points>
<connection>
<GID>350</GID>
<name>clock</name></connection>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-127,199,-123.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-123.5,199,-123.5</points>
<intersection>193 2</intersection>
<intersection>199 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>193,-123.5,193,-74.5</points>
<intersection>-123.5 1</intersection>
<intersection>-74.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>186.5,-74.5,193,-74.5</points>
<connection>
<GID>287</GID>
<name>N_in1</name></connection>
<intersection>193 2</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-129,199,-118.5</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-129,222,-129</points>
<intersection>199 0</intersection>
<intersection>222 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>222,-129,222,-101</points>
<intersection>-129 1</intersection>
<intersection>-101 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-101,224,-101</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>222 2</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-120,199,-110</points>
<connection>
<GID>363</GID>
<name>OUT_0</name></connection>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-120 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-120,221,-120</points>
<intersection>199 0</intersection>
<intersection>221 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>221,-120,221,-100</points>
<intersection>-120 3</intersection>
<intersection>-100 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>221,-100,224,-100</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>221 4</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-104,199,-102</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-103 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>199,-103,220,-103</points>
<intersection>199 0</intersection>
<intersection>220 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>220,-103,220,-99</points>
<intersection>-103 6</intersection>
<intersection>-99 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>220,-99,224,-99</points>
<connection>
<GID>360</GID>
<name>IN_2</name></connection>
<intersection>220 7</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-96,199,-94.5</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>-95.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-95.5,219,-95.5</points>
<intersection>199 0</intersection>
<intersection>219 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>219,-98,219,-95.5</points>
<intersection>-98 5</intersection>
<intersection>-95.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>219,-98,224,-98</points>
<connection>
<GID>360</GID>
<name>IN_3</name></connection>
<intersection>219 4</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-97,220,-88</points>
<intersection>-97 5</intersection>
<intersection>-88 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220,-97,224,-97</points>
<connection>
<GID>360</GID>
<name>IN_4</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>199,-88,220,-88</points>
<intersection>199 8</intersection>
<intersection>220 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>199,-88.5,199,-87</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>-88 6</intersection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-81,199,-79.5</points>
<connection>
<GID>367</GID>
<name>OUT_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>-80.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-80.5,221,-80.5</points>
<intersection>199 0</intersection>
<intersection>221 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>221,-96,221,-80.5</points>
<intersection>-96 5</intersection>
<intersection>-80.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>221,-96,224,-96</points>
<connection>
<GID>360</GID>
<name>IN_5</name></connection>
<intersection>221 4</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-73.5,199,-72</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>-73 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>199,-73,222,-73</points>
<intersection>199 0</intersection>
<intersection>222 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>222,-95,222,-73</points>
<intersection>-95 5</intersection>
<intersection>-73 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>222,-95,224,-95</points>
<connection>
<GID>360</GID>
<name>IN_6</name></connection>
<intersection>222 4</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-290.5,115.5,-288.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-290.5,117,-290.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-66,199,-63.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-63.5,224,-63.5</points>
<intersection>199 0</intersection>
<intersection>224 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>224,-94,224,-63.5</points>
<connection>
<GID>360</GID>
<name>IN_7</name></connection>
<intersection>-63.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-103,227,-103</points>
<connection>
<GID>360</GID>
<name>clock</name></connection>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-92,227,-92</points>
<connection>
<GID>360</GID>
<name>load</name></connection>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-207,191.5,-82.5</points>
<intersection>-207 3</intersection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>186.5,-82.5,191.5,-82.5</points>
<connection>
<GID>289</GID>
<name>N_in1</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>191.5,-207,202.5,-207</points>
<intersection>191.5 0</intersection>
<intersection>202.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>202.5,-207,202.5,-203.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-207 3</intersection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-197.5,202.5,-195</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-196.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-196.5,225.5,-196.5</points>
<intersection>202.5 0</intersection>
<intersection>225.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>225.5,-196.5,225.5,-177.5</points>
<intersection>-196.5 1</intersection>
<intersection>-177.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>225.5,-177.5,227.5,-177.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>225.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-189,202.5,-186.5</points>
<connection>
<GID>377</GID>
<name>OUT_0</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-188 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>202.5,-188,224.5,-188</points>
<intersection>202.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,-188,224.5,-176.5</points>
<intersection>-188 3</intersection>
<intersection>-176.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,-176.5,227.5,-176.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-180.5,202.5,-178.5</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>-179.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>202.5,-179.5,223.5,-179.5</points>
<intersection>202.5 0</intersection>
<intersection>223.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>223.5,-179.5,223.5,-175.5</points>
<intersection>-179.5 6</intersection>
<intersection>-175.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>223.5,-175.5,227.5,-175.5</points>
<connection>
<GID>374</GID>
<name>IN_2</name></connection>
<intersection>223.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-172.5,202.5,-171</points>
<connection>
<GID>379</GID>
<name>OUT_0</name></connection>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-172 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>202.5,-172,222.5,-172</points>
<intersection>202.5 0</intersection>
<intersection>222.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>222.5,-174.5,222.5,-172</points>
<intersection>-174.5 5</intersection>
<intersection>-172 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>222.5,-174.5,227.5,-174.5</points>
<connection>
<GID>374</GID>
<name>IN_3</name></connection>
<intersection>222.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,-173.5,223.5,-164.5</points>
<intersection>-173.5 5</intersection>
<intersection>-164.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>223.5,-173.5,227.5,-173.5</points>
<connection>
<GID>374</GID>
<name>IN_4</name></connection>
<intersection>223.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>202.5,-164.5,223.5,-164.5</points>
<intersection>202.5 8</intersection>
<intersection>223.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>202.5,-165,202.5,-163.5</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-164.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-157.5,202.5,-156</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-157 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>202.5,-157,224.5,-157</points>
<intersection>202.5 0</intersection>
<intersection>224.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>224.5,-172.5,224.5,-157</points>
<intersection>-172.5 5</intersection>
<intersection>-157 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>224.5,-172.5,227.5,-172.5</points>
<connection>
<GID>374</GID>
<name>IN_5</name></connection>
<intersection>224.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-150,202.5,-148.5</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>-149.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>202.5,-149.5,225.5,-149.5</points>
<intersection>202.5 0</intersection>
<intersection>225.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>225.5,-171.5,225.5,-149.5</points>
<intersection>-171.5 5</intersection>
<intersection>-149.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>225.5,-171.5,227.5,-171.5</points>
<connection>
<GID>374</GID>
<name>IN_6</name></connection>
<intersection>225.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-276.5,116.5,-266</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-266,116.5,-266</points>
<connection>
<GID>372</GID>
<name>OUT_7</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-142.5,202.5,-140</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-140,227.5,-140</points>
<intersection>202.5 0</intersection>
<intersection>227.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>227.5,-170.5,227.5,-140</points>
<connection>
<GID>374</GID>
<name>IN_7</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-179.5,230.5,-179.5</points>
<connection>
<GID>374</GID>
<name>clock</name></connection>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-168.5,230.5,-168.5</points>
<connection>
<GID>374</GID>
<name>load</name></connection>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-276.5,107.5,-267</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>-267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-267,107.5,-267</points>
<connection>
<GID>372</GID>
<name>OUT_6</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-276.5,98.5,-268</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>-268 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-268,98.5,-268</points>
<connection>
<GID>372</GID>
<name>OUT_5</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-276.5,89.5,-269</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>-269 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-269,89.5,-269</points>
<connection>
<GID>372</GID>
<name>OUT_4</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-276.5,80,-270</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>-270 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-270,80,-270</points>
<connection>
<GID>372</GID>
<name>OUT_3</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-276.5,71,-271</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-271 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-271,71,-271</points>
<connection>
<GID>372</GID>
<name>OUT_2</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-264,43.5,-264</points>
<connection>
<GID>372</GID>
<name>count_enable</name></connection>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-317,117,-317</points>
<intersection>31.5 39</intersection>
<intersection>53.5 34</intersection>
<intersection>62.5 35</intersection>
<intersection>71.5 36</intersection>
<intersection>81 37</intersection>
<intersection>90 38</intersection>
<intersection>99 33</intersection>
<intersection>108 32</intersection>
<intersection>117 31</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>117,-317,117,-293.5</points>
<connection>
<GID>359</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>108,-317,108,-293.5</points>
<connection>
<GID>286</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>99,-317,99,-293.5</points>
<connection>
<GID>271</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>53.5,-317,53.5,-293.5</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>62.5,-317,62.5,-293.5</points>
<connection>
<GID>207</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>71.5,-317,71.5,-293.5</points>
<connection>
<GID>249</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>81,-317,81,-293.5</points>
<connection>
<GID>263</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>90,-317,90,-293.5</points>
<connection>
<GID>267</GID>
<name>clock</name></connection>
<intersection>-317 1</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>31.5,-372,31.5,-317</points>
<intersection>-372 41</intersection>
<intersection>-340.5 81</intersection>
<intersection>-317 1</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>31.5,-372,118.5,-372</points>
<intersection>31.5 39</intersection>
<intersection>55 74</intersection>
<intersection>64 75</intersection>
<intersection>73 76</intersection>
<intersection>82.5 77</intersection>
<intersection>91.5 78</intersection>
<intersection>100.5 73</intersection>
<intersection>109.5 72</intersection>
<intersection>118.5 71</intersection></hsegment>
<vsegment>
<ID>71</ID>
<points>118.5,-389,118.5,-353</points>
<connection>
<GID>183</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>72</ID>
<points>109.5,-372,109.5,-353</points>
<connection>
<GID>177</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>100.5,-372,100.5,-353</points>
<connection>
<GID>172</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>55,-372,55,-353</points>
<connection>
<GID>146</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>64,-372,64,-353</points>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>73,-372,73,-353</points>
<connection>
<GID>159</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>82.5,-372,82.5,-353</points>
<connection>
<GID>163</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>91.5,-372,91.5,-353</points>
<connection>
<GID>167</GID>
<name>clock</name></connection>
<intersection>-372 41</intersection></vsegment>
<hsegment>
<ID>81</ID>
<points>24,-340.5,31.5,-340.5</points>
<intersection>24 82</intersection>
<intersection>25.5 83</intersection>
<intersection>31.5 39</intersection></hsegment>
<vsegment>
<ID>82</ID>
<points>24,-340.5,24,-339</points>
<connection>
<GID>387</GID>
<name>OUT</name></connection>
<intersection>-340.5 81</intersection></vsegment>
<vsegment>
<ID>83</ID>
<points>25.5,-340.5,25.5,-339</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-340.5 81</intersection></vsegment>
<hsegment>
<ID>126</ID>
<points>118.5,-389,288,-389</points>
<intersection>118.5 71</intersection>
<intersection>174 159</intersection>
<intersection>183 160</intersection>
<intersection>192 161</intersection>
<intersection>201.5 162</intersection>
<intersection>210.5 163</intersection>
<intersection>219.5 158</intersection>
<intersection>228.5 157</intersection>
<intersection>237.5 156</intersection>
<intersection>269.5 164</intersection>
<intersection>288 253</intersection></hsegment>
<vsegment>
<ID>156</ID>
<points>237.5,-389,237.5,-370</points>
<connection>
<GID>434</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>157</ID>
<points>228.5,-389,228.5,-370</points>
<connection>
<GID>430</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>158</ID>
<points>219.5,-389,219.5,-370</points>
<connection>
<GID>426</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>159</ID>
<points>174,-389,174,-370</points>
<connection>
<GID>404</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>160</ID>
<points>183,-389,183,-370</points>
<connection>
<GID>410</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>161</ID>
<points>192,-389,192,-370</points>
<connection>
<GID>414</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>162</ID>
<points>201.5,-389,201.5,-370</points>
<connection>
<GID>418</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>163</ID>
<points>210.5,-389,210.5,-370</points>
<connection>
<GID>422</GID>
<name>clock</name></connection>
<intersection>-389 126</intersection></vsegment>
<vsegment>
<ID>164</ID>
<points>269.5,-389,269.5,-296.5</points>
<intersection>-389 126</intersection>
<intersection>-351.5 262</intersection>
<intersection>-343 261</intersection>
<intersection>-334.5 260</intersection>
<intersection>-326.5 259</intersection>
<intersection>-319 258</intersection>
<intersection>-311.5 257</intersection>
<intersection>-304 256</intersection>
<intersection>-296.5 255</intersection></vsegment>
<vsegment>
<ID>253</ID>
<points>288,-389,288,-331.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>-389 126</intersection></vsegment>
<hsegment>
<ID>255</ID>
<points>263,-296.5,269.5,-296.5</points>
<connection>
<GID>458</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>256</ID>
<points>263,-304,269.5,-304</points>
<connection>
<GID>457</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>257</ID>
<points>263,-311.5,269.5,-311.5</points>
<connection>
<GID>456</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>258</ID>
<points>263,-319,269.5,-319</points>
<connection>
<GID>455</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>259</ID>
<points>263,-326.5,269.5,-326.5</points>
<connection>
<GID>454</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>260</ID>
<points>263,-334.5,269.5,-334.5</points>
<connection>
<GID>453</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>261</ID>
<points>263,-343,269.5,-343</points>
<connection>
<GID>452</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment>
<hsegment>
<ID>262</ID>
<points>263,-351.5,269.5,-351.5</points>
<connection>
<GID>451</GID>
<name>clock</name></connection>
<intersection>269.5 164</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>9.5,-341.5,18,-341.5</points>
<connection>
<GID>386</GID>
<name>CLK</name></connection>
<intersection>18 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>18,-341.5,18,-340</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>-341.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-336,11.5,-336</points>
<connection>
<GID>390</GID>
<name>OUT_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-338,18,-337</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-337 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-337,18,-337</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-338,11.5,-338</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>9 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>9,-343.5,9,-338</points>
<intersection>-343.5 10</intersection>
<intersection>-338 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>9,-343.5,16.5,-343.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>9 9</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-343.5,27.5,-339</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>-343.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-343.5,27.5,-343.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-332,26.5,-332</points>
<connection>
<GID>388</GID>
<name>clock</name></connection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-333,26.5,-332</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>-332 1</intersection></vsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>14.5,-331,14.5,-331</points>
<connection>
<GID>388</GID>
<name>count_enable</name></connection>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-336,7.5,-325</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-325 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-325,23.5,-325</points>
<intersection>7.5 0</intersection>
<intersection>17.5 5</intersection>
<intersection>23.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>23.5,-330,23.5,-325</points>
<connection>
<GID>388</GID>
<name>clear</name></connection>
<intersection>-325 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>17.5,-327,17.5,-325</points>
<connection>
<GID>388</GID>
<name>OUT_3</name></connection>
<intersection>-325 1</intersection></vsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-275,42.5,-275</points>
<connection>
<GID>372</GID>
<name>clock</name></connection>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-155,-516,-154,-516</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<connection>
<GID>392</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-350,127.5,-327.5</points>
<intersection>-350 1</intersection>
<intersection>-327.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-350,127.5,-350</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-327.5,141.5,-327.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-326.5,127.5,-290.5</points>
<intersection>-326.5 1</intersection>
<intersection>-290.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-326.5,141.5,-326.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123,-290.5,127.5,-290.5</points>
<connection>
<GID>359</GID>
<name>OUT_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-152,-516,-151,-516</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<connection>
<GID>439</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-72.5,63,-70.5</points>
<intersection>-72.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-72.5,69,-72.5</points>
<connection>
<GID>350</GID>
<name>IN_7</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-70.5,63,-70.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-73.5,62,-72.5</points>
<intersection>-73.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-72.5,62,-72.5</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,-73.5,69,-73.5</points>
<connection>
<GID>350</GID>
<name>IN_6</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-74.5,69,-74.5</points>
<connection>
<GID>350</GID>
<name>IN_5</name></connection>
<connection>
<GID>395</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-76.5,62,-75.5</points>
<intersection>-76.5 1</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-76.5,62,-76.5</points>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62,-75.5,69,-75.5</points>
<connection>
<GID>350</GID>
<name>IN_4</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-78.5,63,-76.5</points>
<intersection>-78.5 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-76.5,69,-76.5</points>
<connection>
<GID>350</GID>
<name>IN_3</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-78.5,63,-78.5</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-80.5,64,-80.5</points>
<connection>
<GID>398</GID>
<name>OUT_0</name></connection>
<intersection>64 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64,-80.5,64,-77.5</points>
<intersection>-80.5 1</intersection>
<intersection>-77.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64,-77.5,69,-77.5</points>
<connection>
<GID>350</GID>
<name>IN_2</name></connection>
<intersection>64 3</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-84.5,66,-79.5</points>
<intersection>-84.5 2</intersection>
<intersection>-79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-79.5,69,-79.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-84.5,66,-84.5</points>
<connection>
<GID>400</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-82.5,65,-78.5</points>
<intersection>-82.5 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-82.5,65,-82.5</points>
<connection>
<GID>399</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-78.5,69,-78.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-70.5,72,-70.5</points>
<connection>
<GID>350</GID>
<name>load</name></connection>
<connection>
<GID>401</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>179.5,-359,180.5,-359</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<connection>
<GID>405</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>182.5,-359,183.5,-359</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<connection>
<GID>406</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-351,235,-351</points>
<intersection>167.5 3</intersection>
<intersection>180.5 2</intersection>
<intersection>189.5 16</intersection>
<intersection>198.5 17</intersection>
<intersection>208 18</intersection>
<intersection>217 19</intersection>
<intersection>226 20</intersection>
<intersection>235 15</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>180.5,-353,180.5,-351</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>167.5,-362.5,167.5,-351</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>-362.5 22</intersection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>235,-353,235,-351</points>
<connection>
<GID>431</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>189.5,-353,189.5,-351</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>198.5,-353,198.5,-351</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>208,-353,208,-351</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>217,-353,217,-351</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>226,-353,226,-351</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-351 1</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>167,-362.5,167.5,-362.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>167.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>171.5,-352.5,239,-352.5</points>
<connection>
<GID>409</GID>
<name>OUT_0</name></connection>
<intersection>184.5 21</intersection>
<intersection>193.5 13</intersection>
<intersection>202.5 14</intersection>
<intersection>212 15</intersection>
<intersection>221 17</intersection>
<intersection>230 18</intersection>
<intersection>239 19</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>193.5,-353,193.5,-352.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>202.5,-353,202.5,-352.5</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>212,-353,212,-352.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>221,-353,221,-352.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>230,-353,230,-352.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>239,-353,239,-352.5</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>184.5,-353,184.5,-352.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<intersection>-352.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-364.5,177,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-364.5,180,-364.5</points>
<intersection>177 0</intersection>
<intersection>180 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-353,178.5,-353</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>177 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>180,-367,180,-364.5</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>188.5,-359,189.5,-359</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<connection>
<GID>411</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>191.5,-359,192.5,-359</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<connection>
<GID>412</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-364.5,186,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,-364.5,189,-364.5</points>
<intersection>186 0</intersection>
<intersection>189 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>186,-353,187.5,-353</points>
<connection>
<GID>411</GID>
<name>IN_1</name></connection>
<intersection>186 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>189,-367,189,-364.5</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>197.5,-359,198.5,-359</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<connection>
<GID>415</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>200.5,-359,201.5,-359</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195,-364.5,195,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,-364.5,198,-364.5</points>
<intersection>195 0</intersection>
<intersection>198 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,-353,196.5,-353</points>
<connection>
<GID>415</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>198,-367,198,-364.5</points>
<connection>
<GID>414</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>207,-359,208,-359</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<connection>
<GID>419</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>210,-359,211,-359</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<connection>
<GID>420</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-364.5,204.5,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-364.5,207.5,-364.5</points>
<intersection>204.5 0</intersection>
<intersection>207.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204.5,-353,206,-353</points>
<connection>
<GID>419</GID>
<name>IN_1</name></connection>
<intersection>204.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>207.5,-367,207.5,-364.5</points>
<connection>
<GID>418</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>216,-359,217,-359</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<connection>
<GID>423</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>219,-359,220,-359</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<connection>
<GID>424</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-364.5,213.5,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-364.5,216.5,-364.5</points>
<intersection>213.5 0</intersection>
<intersection>216.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213.5,-353,215,-353</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>213.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>216.5,-367,216.5,-364.5</points>
<connection>
<GID>422</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>225,-359,226,-359</points>
<connection>
<GID>429</GID>
<name>IN_1</name></connection>
<connection>
<GID>427</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>228,-359,229,-359</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<connection>
<GID>428</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-364.5,222.5,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-364.5,225.5,-364.5</points>
<intersection>222.5 0</intersection>
<intersection>225.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222.5,-353,224,-353</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>222.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>225.5,-367,225.5,-364.5</points>
<connection>
<GID>426</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>234,-359,235,-359</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<connection>
<GID>431</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>237,-359,238,-359</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<connection>
<GID>432</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-364.5,231.5,-353</points>
<intersection>-364.5 1</intersection>
<intersection>-353 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,-364.5,234.5,-364.5</points>
<intersection>231.5 0</intersection>
<intersection>234.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>231.5,-353,233,-353</points>
<connection>
<GID>431</GID>
<name>IN_1</name></connection>
<intersection>231.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>234.5,-367,234.5,-364.5</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<intersection>-364.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-367,174,-349.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>-349.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>168,-349.5,174,-349.5</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,-353,182.5,-348.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<intersection>-348.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-348.5,182.5,-348.5</points>
<connection>
<GID>436</GID>
<name>OUT_1</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-367,181.5,-365</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-367,183,-367</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-367,199.5,-365</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-367,201.5,-367</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>199.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-367,190.5,-365</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,-367,192,-367</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>190.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-367,209,-365</points>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,-367,210.5,-367</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>209 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-367,218,-365</points>
<connection>
<GID>425</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-367,219.5,-367</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-367,227,-365</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-367,228.5,-367</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-367,236,-365</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>-367 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-367,237.5,-367</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>236 0</intersection></hsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,-353,237,-342.5</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-342.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-342.5,237,-342.5</points>
<connection>
<GID>436</GID>
<name>OUT_7</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-353,228,-343.5</points>
<connection>
<GID>428</GID>
<name>IN_1</name></connection>
<intersection>-343.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-343.5,228,-343.5</points>
<connection>
<GID>436</GID>
<name>OUT_6</name></connection>
<intersection>228 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-353,219,-344.5</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-344.5,219,-344.5</points>
<connection>
<GID>436</GID>
<name>OUT_5</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-353,210,-345.5</points>
<connection>
<GID>420</GID>
<name>IN_1</name></connection>
<intersection>-345.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-345.5,210,-345.5</points>
<connection>
<GID>436</GID>
<name>OUT_4</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,-353,200.5,-346.5</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>-346.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-346.5,200.5,-346.5</points>
<connection>
<GID>436</GID>
<name>OUT_3</name></connection>
<intersection>200.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-353,191.5,-347.5</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>-347.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-347.5,191.5,-347.5</points>
<connection>
<GID>436</GID>
<name>OUT_2</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-157.5,-521.5,-157.5,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-157.5,-521.5,-154.5,-521.5</points>
<intersection>-157.5 0</intersection>
<intersection>-154.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-157.5,-510,-156,-510</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>-157.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-154.5,-524,-154.5,-521.5</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-351.5,163,-351.5</points>
<connection>
<GID>436</GID>
<name>clock</name></connection>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-146,-516,-145,-516</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<connection>
<GID>459</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-353,159,-349.5</points>
<intersection>-353 2</intersection>
<intersection>-349.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159,-349.5,160,-349.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-353,159,-353</points>
<connection>
<GID>447</GID>
<name>OUT_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-351,157.5,-348.5</points>
<intersection>-351 1</intersection>
<intersection>-348.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-351,157.5,-351</points>
<connection>
<GID>446</GID>
<name>OUT_0</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-348.5,160,-348.5</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-349,157,-347.5</points>
<intersection>-349 2</intersection>
<intersection>-347.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-347.5,160,-347.5</points>
<connection>
<GID>436</GID>
<name>IN_2</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-349,157,-349</points>
<connection>
<GID>445</GID>
<name>OUT_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-347,156,-346.5</points>
<intersection>-347 1</intersection>
<intersection>-346.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-347,156,-347</points>
<connection>
<GID>444</GID>
<name>OUT_0</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-346.5,160,-346.5</points>
<connection>
<GID>436</GID>
<name>IN_3</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156,-345.5,156,-345</points>
<intersection>-345.5 1</intersection>
<intersection>-345 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156,-345.5,160,-345.5</points>
<connection>
<GID>436</GID>
<name>IN_4</name></connection>
<intersection>156 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-345,156,-345</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<intersection>156 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-343.5,158,-341</points>
<intersection>-343.5 1</intersection>
<intersection>-341 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,-343.5,160,-343.5</points>
<connection>
<GID>436</GID>
<name>IN_6</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-341,158,-341</points>
<connection>
<GID>441</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-344.5,157,-343</points>
<intersection>-344.5 2</intersection>
<intersection>-343 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-343,157,-343</points>
<connection>
<GID>442</GID>
<name>OUT_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,-344.5,160,-344.5</points>
<connection>
<GID>436</GID>
<name>IN_5</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-342.5,159,-339</points>
<intersection>-342.5 2</intersection>
<intersection>-339 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-339,159,-339</points>
<connection>
<GID>440</GID>
<name>OUT_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>159,-342.5,160,-342.5</points>
<connection>
<GID>436</GID>
<name>IN_7</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-340.5,163,-340.5</points>
<connection>
<GID>436</GID>
<name>load</name></connection>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-353.5,260,-351.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>-353.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248.5,-353.5,260,-353.5</points>
<intersection>248.5 2</intersection>
<intersection>260 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>248.5,-353.5,248.5,-328.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>-353.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-345.5,260,-343</points>
<connection>
<GID>451</GID>
<name>OUT_0</name></connection>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>-344.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-344.5,283,-344.5</points>
<intersection>260 0</intersection>
<intersection>283 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283,-344.5,283,-325.5</points>
<intersection>-344.5 1</intersection>
<intersection>-325.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>283,-325.5,285,-325.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<intersection>283 2</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-337,260,-334.5</points>
<connection>
<GID>452</GID>
<name>OUT_0</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>-336 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>260,-336,282,-336</points>
<intersection>260 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-336,282,-324.5</points>
<intersection>-336 3</intersection>
<intersection>-324.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,-324.5,285,-324.5</points>
<connection>
<GID>449</GID>
<name>IN_1</name></connection>
<intersection>282 4</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-328.5,260,-326.5</points>
<connection>
<GID>453</GID>
<name>OUT_0</name></connection>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-327.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>260,-327.5,281,-327.5</points>
<intersection>260 0</intersection>
<intersection>281 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>281,-327.5,281,-323.5</points>
<intersection>-327.5 6</intersection>
<intersection>-323.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>281,-323.5,285,-323.5</points>
<connection>
<GID>449</GID>
<name>IN_2</name></connection>
<intersection>281 7</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-320.5,260,-319</points>
<connection>
<GID>454</GID>
<name>OUT_0</name></connection>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>-320 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>260,-320,280,-320</points>
<intersection>260 0</intersection>
<intersection>280 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>280,-322.5,280,-320</points>
<intersection>-322.5 5</intersection>
<intersection>-320 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>280,-322.5,285,-322.5</points>
<connection>
<GID>449</GID>
<name>IN_3</name></connection>
<intersection>280 4</intersection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-321.5,281,-312.5</points>
<intersection>-321.5 5</intersection>
<intersection>-312.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>281,-321.5,285,-321.5</points>
<connection>
<GID>449</GID>
<name>IN_4</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>260,-312.5,281,-312.5</points>
<intersection>260 8</intersection>
<intersection>281 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>260,-313,260,-311.5</points>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<intersection>-312.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-305.5,260,-304</points>
<connection>
<GID>456</GID>
<name>OUT_0</name></connection>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>-305 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>260,-305,282,-305</points>
<intersection>260 0</intersection>
<intersection>282 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>282,-320.5,282,-305</points>
<intersection>-320.5 5</intersection>
<intersection>-305 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>282,-320.5,285,-320.5</points>
<connection>
<GID>449</GID>
<name>IN_5</name></connection>
<intersection>282 4</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-298,260,-296.5</points>
<connection>
<GID>457</GID>
<name>OUT_0</name></connection>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>-297.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>260,-297.5,283,-297.5</points>
<intersection>260 0</intersection>
<intersection>283 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>283,-319.5,283,-297.5</points>
<intersection>-319.5 5</intersection>
<intersection>-297.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>283,-319.5,285,-319.5</points>
<connection>
<GID>449</GID>
<name>IN_6</name></connection>
<intersection>283 4</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-143,-516,-142,-516</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<connection>
<GID>461</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,-290.5,260,-288</points>
<connection>
<GID>458</GID>
<name>OUT_0</name></connection>
<intersection>-288 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>260,-288,285,-288</points>
<intersection>260 0</intersection>
<intersection>285 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>285,-318.5,285,-288</points>
<connection>
<GID>449</GID>
<name>IN_7</name></connection>
<intersection>-288 1</intersection></vsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148.5,-521.5,-148.5,-510</points>
<intersection>-521.5 1</intersection>
<intersection>-510 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-148.5,-521.5,-145.5,-521.5</points>
<intersection>-148.5 0</intersection>
<intersection>-145.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-148.5,-510,-147,-510</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<intersection>-148.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-145.5,-524,-145.5,-521.5</points>
<connection>
<GID>450</GID>
<name>OUT_0</name></connection>
<intersection>-521.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-316.5,288,-316.5</points>
<connection>
<GID>449</GID>
<name>load</name></connection>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-367,244.5,-329.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-367 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>243.5,-367,244.5,-367</points>
<connection>
<GID>434</GID>
<name>OUT_0</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-208.5,-524,-208.5,-506.5</points>
<intersection>-524 4</intersection>
<intersection>-506.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-212,-506.5,-208.5,-506.5</points>
<connection>
<GID>467</GID>
<name>OUT_0</name></connection>
<intersection>-208.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-208.5,-524,-206,-524</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-327.5,288,-327.5</points>
<connection>
<GID>449</GID>
<name>clock</name></connection>
<connection>
<GID>463</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197.5,-510,-197.5,-505.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>-505.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-505.5,-197.5,-505.5</points>
<connection>
<GID>467</GID>
<name>OUT_1</name></connection>
<intersection>-197.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198.5,-524,-198.5,-522</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-198.5,-524,-197,-524</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-180.5,-524,-180.5,-522</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-180.5,-524,-178.5,-524</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-189.5,-524,-189.5,-522</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-189.5,-524,-188,-524</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-171,-524,-171,-522</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-171,-524,-169.5,-524</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-171 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-162,-524,-162,-522</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-162,-524,-160.5,-524</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-162 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153,-524,-153,-522</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-153,-524,-151.5,-524</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>-153 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-144,-524,-144,-522</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-144,-524,-142.5,-524</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>-144 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-143,-510,-143,-499.5</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>-499.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-499.5,-143,-499.5</points>
<connection>
<GID>467</GID>
<name>OUT_7</name></connection>
<intersection>-143 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-152,-510,-152,-500.5</points>
<connection>
<GID>439</GID>
<name>IN_1</name></connection>
<intersection>-500.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-500.5,-152,-500.5</points>
<connection>
<GID>467</GID>
<name>OUT_6</name></connection>
<intersection>-152 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-161,-510,-161,-501.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>-501.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-501.5,-161,-501.5</points>
<connection>
<GID>467</GID>
<name>OUT_5</name></connection>
<intersection>-161 0</intersection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-170,-510,-170,-502.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>-502.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-502.5,-170,-502.5</points>
<connection>
<GID>467</GID>
<name>OUT_4</name></connection>
<intersection>-170 0</intersection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-179.5,-510,-179.5,-503.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-503.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-503.5,-179.5,-503.5</points>
<connection>
<GID>467</GID>
<name>OUT_3</name></connection>
<intersection>-179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-188.5,-510,-188.5,-504.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-504.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212,-504.5,-188.5,-504.5</points>
<connection>
<GID>467</GID>
<name>OUT_2</name></connection>
<intersection>-188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<hsegment>
<ID>58</ID>
<points>-188.5,-571,-24,-571</points>
<intersection>-188.5 1038</intersection>
<intersection>-24 148</intersection></hsegment>
<hsegment>
<ID>110</ID>
<points>-24,-575,62,-575</points>
<intersection>-24 148</intersection>
<intersection>-1.5 1011</intersection>
<intersection>7.5 1012</intersection>
<intersection>16.5 1013</intersection>
<intersection>26 1014</intersection>
<intersection>35 1015</intersection>
<intersection>44 1016</intersection>
<intersection>53 1017</intersection>
<intersection>62 1018</intersection></hsegment>
<vsegment>
<ID>148</ID>
<points>-24,-630,-24,-571</points>
<intersection>-630 150</intersection>
<intersection>-575 110</intersection>
<intersection>-571 58</intersection></vsegment>
<hsegment>
<ID>150</ID>
<points>-24,-630,63.5,-630</points>
<intersection>-24 148</intersection>
<intersection>0 1019</intersection>
<intersection>9 1020</intersection>
<intersection>18 1021</intersection>
<intersection>27.5 1022</intersection>
<intersection>36.5 1023</intersection>
<intersection>45.5 1024</intersection>
<intersection>54.5 1025</intersection>
<intersection>63.5 180</intersection></hsegment>
<vsegment>
<ID>180</ID>
<points>63.5,-651,63.5,-612.5</points>
<connection>
<GID>549</GID>
<name>clock</name></connection>
<intersection>-651 235</intersection>
<intersection>-630 150</intersection></vsegment>
<hsegment>
<ID>235</ID>
<points>63.5,-651,212,-651</points>
<intersection>63.5 180</intersection>
<intersection>212 1040</intersection></hsegment>
<vsegment>
<ID>1011</ID>
<points>-1.5,-575,-1.5,-553</points>
<connection>
<GID>554</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1012</ID>
<points>7.5,-575,7.5,-553</points>
<connection>
<GID>562</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1013</ID>
<points>16.5,-575,16.5,-553</points>
<connection>
<GID>567</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1014</ID>
<points>26,-575,26,-553</points>
<connection>
<GID>571</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1015</ID>
<points>35,-575,35,-553</points>
<connection>
<GID>575</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1016</ID>
<points>44,-575,44,-553</points>
<connection>
<GID>579</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1017</ID>
<points>53,-575,53,-553</points>
<connection>
<GID>583</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1018</ID>
<points>62,-575,62,-553</points>
<connection>
<GID>587</GID>
<name>clock</name></connection>
<intersection>-575 110</intersection></vsegment>
<vsegment>
<ID>1019</ID>
<points>0,-630,0,-612.5</points>
<connection>
<GID>519</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1020</ID>
<points>9,-630,9,-612.5</points>
<connection>
<GID>525</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1021</ID>
<points>18,-630,18,-612.5</points>
<connection>
<GID>529</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1022</ID>
<points>27.5,-630,27.5,-612.5</points>
<connection>
<GID>533</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1023</ID>
<points>36.5,-630,36.5,-612.5</points>
<connection>
<GID>537</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1024</ID>
<points>45.5,-630,45.5,-612.5</points>
<connection>
<GID>541</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1025</ID>
<points>54.5,-630,54.5,-612.5</points>
<connection>
<GID>545</GID>
<name>clock</name></connection>
<intersection>-630 150</intersection></vsegment>
<vsegment>
<ID>1038</ID>
<points>-188.5,-571,-188.5,-557</points>
<intersection>-571 58</intersection>
<intersection>-557 1039</intersection></vsegment>
<hsegment>
<ID>1039</ID>
<points>-203.5,-557,-188.5,-557</points>
<connection>
<GID>510</GID>
<name>OUT</name></connection>
<intersection>-188.5 1038</intersection></hsegment>
<vsegment>
<ID>1040</ID>
<points>212,-651,212,-624</points>
<intersection>-651 235</intersection>
<intersection>-624 1041</intersection></vsegment>
<hsegment>
<ID>1041</ID>
<points>212,-624,215.5,-624</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>212 1040</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-232,-548.5,-229.5,-548.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>-232 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-232,-550,-232,-548.5</points>
<intersection>-550 12</intersection>
<intersection>-548.5 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-238,-550,-232,-550</points>
<connection>
<GID>469</GID>
<name>CLK</name></connection>
<intersection>-232 11</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-236,-544.5,-236,-544.5</points>
<connection>
<GID>473</GID>
<name>OUT_0</name></connection>
<connection>
<GID>474</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-229.5,-546.5,-229.5,-545.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>-545.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-230,-545.5,-229.5,-545.5</points>
<connection>
<GID>474</GID>
<name>OUT</name></connection>
<intersection>-229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-243.5,-546.5,-236,-546.5</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>-243.5 14</intersection>
<intersection>-237.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-237.5,-552,-237.5,-546.5</points>
<intersection>-552 16</intersection>
<intersection>-546.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-243.5,-546.5,-243.5,-541</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>-546.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-237.5,-552,-231,-552</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-237.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220,-552,-220,-547.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-552 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227,-552,-220,-552</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-220 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-224,-540.5,-221,-540.5</points>
<connection>
<GID>471</GID>
<name>clock</name></connection>
<intersection>-221 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-221,-541.5,-221,-540.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-540.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-233,-539.5,-233,-539.5</points>
<connection>
<GID>471</GID>
<name>count_enable</name></connection>
<connection>
<GID>472</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-240,-544.5,-240,-528.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>-528.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-240,-528.5,-224,-528.5</points>
<intersection>-240 0</intersection>
<intersection>-228.5 3</intersection>
<intersection>-224 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-224,-538.5,-224,-528.5</points>
<connection>
<GID>471</GID>
<name>clear</name></connection>
<intersection>-528.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-228.5,-529,-228.5,-528.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-528.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,-535.5,-230,-535</points>
<connection>
<GID>471</GID>
<name>OUT_3</name></connection>
<intersection>-535 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-230,-535,-229.5,-535</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-230 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79.5,-558,-65,-558</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>-79.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-79.5,-558,-79.5,-502.5</points>
<intersection>-558 1</intersection>
<intersection>-502.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-98,-502.5,-79.5,-502.5</points>
<connection>
<GID>45</GID>
<name>N_in1</name></connection>
<intersection>-79.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-552,-65,-549.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<connection>
<GID>476</GID>
<name>OUT_0</name></connection>
<intersection>-551 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-551,-42,-551</points>
<intersection>-65 0</intersection>
<intersection>-42 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-42,-551,-42,-532</points>
<intersection>-551 1</intersection>
<intersection>-532 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-42,-532,-40,-532</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>-42 2</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-543.5,-65,-541</points>
<connection>
<GID>477</GID>
<name>OUT_0</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>-542 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-65,-542,-43,-542</points>
<intersection>-65 0</intersection>
<intersection>-43 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-43,-542,-43,-531</points>
<intersection>-542 3</intersection>
<intersection>-531 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-43,-531,-40,-531</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>-43 4</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-535,-65,-533</points>
<connection>
<GID>478</GID>
<name>OUT_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>-534 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-65,-534,-44,-534</points>
<intersection>-65 0</intersection>
<intersection>-44 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-44,-534,-44,-530</points>
<intersection>-534 6</intersection>
<intersection>-530 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-44,-530,-40,-530</points>
<connection>
<GID>475</GID>
<name>IN_2</name></connection>
<intersection>-44 7</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-527,-65,-525.5</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-65,-526.5,-45,-526.5</points>
<intersection>-65 0</intersection>
<intersection>-45 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-45,-529,-45,-526.5</points>
<intersection>-529 5</intersection>
<intersection>-526.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-45,-529,-40,-529</points>
<connection>
<GID>475</GID>
<name>IN_3</name></connection>
<intersection>-45 4</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-528,-44,-518.5</points>
<intersection>-528 5</intersection>
<intersection>-518.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-44,-528,-40,-528</points>
<connection>
<GID>475</GID>
<name>IN_4</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-65,-518.5,-44,-518.5</points>
<intersection>-65 8</intersection>
<intersection>-44 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-65,-519.5,-65,-518</points>
<connection>
<GID>480</GID>
<name>OUT_0</name></connection>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>-518.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-512,-65,-510.5</points>
<connection>
<GID>481</GID>
<name>OUT_0</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>-511.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-65,-511.5,-43,-511.5</points>
<intersection>-65 0</intersection>
<intersection>-43 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-43,-527,-43,-511.5</points>
<intersection>-527 5</intersection>
<intersection>-511.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-43,-527,-40,-527</points>
<connection>
<GID>475</GID>
<name>IN_5</name></connection>
<intersection>-43 4</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-504.5,-65,-503</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>-504 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-65,-504,-42,-504</points>
<intersection>-65 0</intersection>
<intersection>-42 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-42,-526,-42,-504</points>
<intersection>-526 5</intersection>
<intersection>-504 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-42,-526,-40,-526</points>
<connection>
<GID>475</GID>
<name>IN_6</name></connection>
<intersection>-42 4</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,-497,-65,-496.5</points>
<connection>
<GID>483</GID>
<name>OUT_0</name></connection>
<intersection>-496.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-496.5,-40,-496.5</points>
<intersection>-65 0</intersection>
<intersection>-40 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-40,-525,-40,-496.5</points>
<connection>
<GID>475</GID>
<name>IN_7</name></connection>
<intersection>-496.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-523,-37,-523</points>
<connection>
<GID>475</GID>
<name>load</name></connection>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-82.5,-642,-82.5,-510.5</points>
<intersection>-642 3</intersection>
<intersection>-510.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-98,-510.5,-82.5,-510.5</points>
<connection>
<GID>54</GID>
<name>N_in1</name></connection>
<intersection>-82.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-82.5,-642,-63,-642</points>
<intersection>-82.5 0</intersection>
<intersection>-63 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-63,-642,-63,-641</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>-642 3</intersection></vsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-635,-63,-632.5</points>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-634 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-634,-40,-634</points>
<intersection>-63 0</intersection>
<intersection>-40 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-40,-634,-40,-615</points>
<intersection>-634 1</intersection>
<intersection>-615 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-40,-615,-38,-615</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>-40 2</intersection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-626.5,-63,-624</points>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>-625.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-63,-625.5,-41,-625.5</points>
<intersection>-63 0</intersection>
<intersection>-41 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-41,-625.5,-41,-614</points>
<intersection>-625.5 3</intersection>
<intersection>-614 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-41,-614,-38,-614</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>-41 4</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-618,-63,-616</points>
<connection>
<GID>489</GID>
<name>OUT_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>-617 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-63,-617,-42,-617</points>
<intersection>-63 0</intersection>
<intersection>-42 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-42,-617,-42,-613</points>
<intersection>-617 6</intersection>
<intersection>-613 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-42,-613,-38,-613</points>
<connection>
<GID>486</GID>
<name>IN_2</name></connection>
<intersection>-42 7</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-610,-63,-608.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection>
<intersection>-609.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-63,-609.5,-43,-609.5</points>
<intersection>-63 0</intersection>
<intersection>-43 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-43,-612,-43,-609.5</points>
<intersection>-612 5</intersection>
<intersection>-609.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-43,-612,-38,-612</points>
<connection>
<GID>486</GID>
<name>IN_3</name></connection>
<intersection>-43 4</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-611,-42,-602</points>
<intersection>-611 5</intersection>
<intersection>-602 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-42,-611,-38,-611</points>
<connection>
<GID>486</GID>
<name>IN_4</name></connection>
<intersection>-42 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-63,-602,-42,-602</points>
<intersection>-63 8</intersection>
<intersection>-42 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-63,-602.5,-63,-601</points>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>-602 6</intersection></vsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-595,-63,-593.5</points>
<connection>
<GID>492</GID>
<name>OUT_0</name></connection>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-594.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-63,-594.5,-41,-594.5</points>
<intersection>-63 0</intersection>
<intersection>-41 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-41,-610,-41,-594.5</points>
<intersection>-610 5</intersection>
<intersection>-594.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-41,-610,-38,-610</points>
<connection>
<GID>486</GID>
<name>IN_5</name></connection>
<intersection>-41 4</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-587.5,-63,-586</points>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-587 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-63,-587,-40,-587</points>
<intersection>-63 0</intersection>
<intersection>-40 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-40,-609,-40,-587</points>
<intersection>-609 5</intersection>
<intersection>-587 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-40,-609,-38,-609</points>
<connection>
<GID>486</GID>
<name>IN_6</name></connection>
<intersection>-40 4</intersection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-580,-63,-577.5</points>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>-577.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,-577.5,-38,-577.5</points>
<intersection>-63 0</intersection>
<intersection>-38 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-38,-608,-38,-577.5</points>
<connection>
<GID>486</GID>
<name>IN_7</name></connection>
<intersection>-577.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-228,-527.5,-212.5,-527.5</points>
<intersection>-228 7</intersection>
<intersection>-212.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-212.5,-544.5,-212.5,-527.5</points>
<intersection>-544.5 5</intersection>
<intersection>-527.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-212.5,-544.5,-200,-544.5</points>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<intersection>-212.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-228,-527.5,-228,-525</points>
<intersection>-527.5 1</intersection>
<intersection>-525 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-230,-525,-227,-525</points>
<connection>
<GID>697</GID>
<name>OUT</name></connection>
<connection>
<GID>495</GID>
<name>IN_1</name></connection>
<intersection>-228 7</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,-606,-35,-606</points>
<connection>
<GID>486</GID>
<name>load</name></connection>
<connection>
<GID>496</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-226,-499.5,-226,-497.5</points>
<intersection>-499.5 1</intersection>
<intersection>-497.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-226,-499.5,-220,-499.5</points>
<connection>
<GID>467</GID>
<name>IN_7</name></connection>
<intersection>-226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233,-497.5,-226,-497.5</points>
<connection>
<GID>497</GID>
<name>OUT_0</name></connection>
<intersection>-226 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227,-500.5,-227,-499.5</points>
<intersection>-500.5 2</intersection>
<intersection>-499.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233,-499.5,-227,-499.5</points>
<connection>
<GID>498</GID>
<name>OUT_0</name></connection>
<intersection>-227 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-227,-500.5,-220,-500.5</points>
<connection>
<GID>467</GID>
<name>IN_6</name></connection>
<intersection>-227 0</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-233,-501.5,-220,-501.5</points>
<connection>
<GID>467</GID>
<name>IN_5</name></connection>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227.5,-503.5,-227.5,-502.5</points>
<intersection>-503.5 1</intersection>
<intersection>-502.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233,-503.5,-227.5,-503.5</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<intersection>-227.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-227.5,-502.5,-220,-502.5</points>
<connection>
<GID>467</GID>
<name>IN_4</name></connection>
<intersection>-227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-226.5,-505.5,-226.5,-503.5</points>
<intersection>-505.5 2</intersection>
<intersection>-503.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-226.5,-503.5,-220,-503.5</points>
<connection>
<GID>467</GID>
<name>IN_3</name></connection>
<intersection>-226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233,-505.5,-226.5,-505.5</points>
<connection>
<GID>501</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-233,-507.5,-225.5,-507.5</points>
<connection>
<GID>502</GID>
<name>OUT_0</name></connection>
<intersection>-225.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-225.5,-507.5,-225.5,-504.5</points>
<intersection>-507.5 1</intersection>
<intersection>-504.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-225.5,-504.5,-220,-504.5</points>
<connection>
<GID>467</GID>
<name>IN_2</name></connection>
<intersection>-225.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-223.5,-511.5,-223.5,-506.5</points>
<intersection>-511.5 2</intersection>
<intersection>-506.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-223.5,-506.5,-220,-506.5</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>-223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233,-511.5,-223.5,-511.5</points>
<connection>
<GID>504</GID>
<name>OUT_0</name></connection>
<intersection>-223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224.5,-509.5,-224.5,-505.5</points>
<intersection>-509.5 1</intersection>
<intersection>-505.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233,-509.5,-224.5,-509.5</points>
<connection>
<GID>503</GID>
<name>OUT_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-224.5,-505.5,-220,-505.5</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<intersection>-224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-217,-497.5,-217,-497.5</points>
<connection>
<GID>467</GID>
<name>load</name></connection>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-227,-535.5,-227,-535</points>
<connection>
<GID>471</GID>
<name>OUT_0</name></connection>
<intersection>-535 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-227.5,-535,-227,-535</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-227 0</intersection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-221,-524,-221,-516.5</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<connection>
<GID>698</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92.5,-580,206.5,-580</points>
<connection>
<GID>515</GID>
<name>IN_1</name></connection>
<intersection>92.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>92.5,-583.5,92.5,-580</points>
<intersection>-583.5 7</intersection>
<intersection>-580 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>87,-583.5,92.5,-583.5</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>92.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-210,-556,-210,-550</points>
<intersection>-556 7</intersection>
<intersection>-550 5</intersection>
<intersection>-550 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-211.5,-550,-209.5,-550</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>-210 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-210,-556,-209.5,-556</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>-210 1</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>5.5,-601.5,6.5,-601.5</points>
<connection>
<GID>522</GID>
<name>IN_1</name></connection>
<connection>
<GID>520</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>8.5,-601.5,9.5,-601.5</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<connection>
<GID>521</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230.5,-523,-230.5,-482.5</points>
<intersection>-523 10</intersection>
<intersection>-520 5</intersection>
<intersection>-516.5 13</intersection>
<intersection>-482.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,-482.5,-230.5,-482.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-230.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-230.5,-520,-209.5,-520</points>
<intersection>-230.5 0</intersection>
<intersection>-209.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-209.5,-548,-209.5,-520</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>-520 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-230.5,-523,-227,-523</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>-230.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-232.5,-516.5,-230.5,-516.5</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<intersection>-230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-243.5,-517.5,-238.5,-517.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-607,3,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-607,6,-607</points>
<intersection>3 0</intersection>
<intersection>6 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-595.5,4.5,-595.5</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6,-609.5,6,-607</points>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>14.5,-601.5,15.5,-601.5</points>
<connection>
<GID>528</GID>
<name>IN_1</name></connection>
<connection>
<GID>526</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>17.5,-601.5,18.5,-601.5</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<connection>
<GID>527</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-607,12,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-607,15,-607</points>
<intersection>12 0</intersection>
<intersection>15 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-595.5,13.5,-595.5</points>
<connection>
<GID>526</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-609.5,15,-607</points>
<connection>
<GID>525</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>23.5,-601.5,24.5,-601.5</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<connection>
<GID>530</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26.5,-601.5,27.5,-601.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-607,21,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-607,24,-607</points>
<intersection>21 0</intersection>
<intersection>24 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-595.5,22.5,-595.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-609.5,24,-607</points>
<connection>
<GID>529</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>33,-601.5,34,-601.5</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<connection>
<GID>534</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>36,-601.5,37,-601.5</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<connection>
<GID>535</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-607,30.5,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-607,33.5,-607</points>
<intersection>30.5 0</intersection>
<intersection>33.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-595.5,32,-595.5</points>
<connection>
<GID>534</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-609.5,33.5,-607</points>
<connection>
<GID>533</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>42,-601.5,43,-601.5</points>
<connection>
<GID>540</GID>
<name>IN_1</name></connection>
<connection>
<GID>538</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45,-601.5,46,-601.5</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<connection>
<GID>539</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-607,39.5,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-607,42.5,-607</points>
<intersection>39.5 0</intersection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-595.5,41,-595.5</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-609.5,42.5,-607</points>
<connection>
<GID>537</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>51,-601.5,52,-601.5</points>
<connection>
<GID>544</GID>
<name>IN_1</name></connection>
<connection>
<GID>542</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>54,-601.5,55,-601.5</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<connection>
<GID>543</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-607,48.5,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48.5,-607,51.5,-607</points>
<intersection>48.5 0</intersection>
<intersection>51.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-595.5,50,-595.5</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>48.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51.5,-609.5,51.5,-607</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>60,-601.5,61,-601.5</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<connection>
<GID>546</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>63,-601.5,64,-601.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<connection>
<GID>547</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-607,57.5,-595.5</points>
<intersection>-607 1</intersection>
<intersection>-595.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-607,60.5,-607</points>
<intersection>57.5 0</intersection>
<intersection>60.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-595.5,59,-595.5</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>57.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-609.5,60.5,-607</points>
<connection>
<GID>545</GID>
<name>OUT_0</name></connection>
<intersection>-607 1</intersection></vsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-223.5,-547.5,-217.5,-547.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<intersection>-217.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-217.5,-551,-217.5,-547.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>-547.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-206.5,-534.5,-206.5,-527</points>
<intersection>-534.5 1</intersection>
<intersection>-527 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-206.5,-534.5,-142.5,-534.5</points>
<intersection>-206.5 0</intersection>
<intersection>-203.5 3</intersection>
<intersection>-197 10</intersection>
<intersection>-188 9</intersection>
<intersection>-178.5 8</intersection>
<intersection>-169.5 7</intersection>
<intersection>-160.5 6</intersection>
<intersection>-151.5 5</intersection>
<intersection>-142.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-206.5,-527,-206,-527</points>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<intersection>-206.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-203.5,-549,-203.5,-534.5</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-142.5,-565.5,-142.5,-527</points>
<connection>
<GID>465</GID>
<name>clock</name></connection>
<intersection>-565.5 12</intersection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-151.5,-534.5,-151.5,-527</points>
<connection>
<GID>450</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-160.5,-534.5,-160.5,-527</points>
<connection>
<GID>352</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-169.5,-534.5,-169.5,-527</points>
<connection>
<GID>192</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-178.5,-534.5,-178.5,-527</points>
<connection>
<GID>152</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-188,-534.5,-188,-527</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-197,-534.5,-197,-527</points>
<connection>
<GID>114</GID>
<name>clock</name></connection>
<intersection>-534.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-142.5,-565.5,-57,-565.5</points>
<intersection>-142.5 4</intersection>
<intersection>-57 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>-57,-641,-57,-503</points>
<intersection>-641 24</intersection>
<intersection>-632.5 31</intersection>
<intersection>-624 30</intersection>
<intersection>-616 29</intersection>
<intersection>-608.5 28</intersection>
<intersection>-601 27</intersection>
<intersection>-593.5 26</intersection>
<intersection>-586 25</intersection>
<intersection>-565.5 12</intersection>
<intersection>-558 16</intersection>
<intersection>-549.5 22</intersection>
<intersection>-541 21</intersection>
<intersection>-533 20</intersection>
<intersection>-525.5 19</intersection>
<intersection>-518 18</intersection>
<intersection>-510.5 17</intersection>
<intersection>-503 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-62,-503,-57,-503</points>
<connection>
<GID>483</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-62,-558,-37,-558</points>
<connection>
<GID>476</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection>
<intersection>-37 35</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-62,-510.5,-57,-510.5</points>
<connection>
<GID>482</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-62,-518,-57,-518</points>
<connection>
<GID>481</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>-62,-525.5,-57,-525.5</points>
<connection>
<GID>480</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-62,-533,-57,-533</points>
<connection>
<GID>479</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-62,-541,-57,-541</points>
<connection>
<GID>478</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-62,-549.5,-57,-549.5</points>
<connection>
<GID>477</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-60,-641,-35,-641</points>
<connection>
<GID>487</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection>
<intersection>-35 33</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-60,-586,-57,-586</points>
<connection>
<GID>494</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-60,-593.5,-57,-593.5</points>
<connection>
<GID>493</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-60,-601,-57,-601</points>
<connection>
<GID>492</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-60,-608.5,-57,-608.5</points>
<connection>
<GID>491</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-60,-616,-57,-616</points>
<connection>
<GID>490</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-60,-624,-57,-624</points>
<connection>
<GID>489</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>-60,-632.5,-57,-632.5</points>
<connection>
<GID>488</GID>
<name>clock</name></connection>
<intersection>-57 13</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>-35,-641,-35,-621</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<intersection>-641 24</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-37,-558,-37,-538</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>-558 16</intersection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-609.5,7.5,-607.5</points>
<connection>
<GID>522</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-609.5,9,-609.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-609.5,25.5,-607.5</points>
<connection>
<GID>532</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-609.5,27.5,-609.5</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-609.5,16.5,-607.5</points>
<connection>
<GID>528</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-609.5,18,-609.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-609.5,35,-607.5</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-609.5,36.5,-609.5</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-609.5,44,-607.5</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-609.5,45.5,-609.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-609.5,53,-607.5</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-609.5,54.5,-609.5</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-609.5,62,-607.5</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<intersection>-609.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-609.5,63.5,-609.5</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-183.5,-544.5,-183.5,-540</points>
<intersection>-544.5 16</intersection>
<intersection>-543.5 8</intersection>
<intersection>-542.5 7</intersection>
<intersection>-540 18</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-183.5,-542.5,-182.5,-542.5</points>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>-183.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-184,-543.5,-183.5,-543.5</points>
<connection>
<GID>524</GID>
<name>OUT_0</name></connection>
<intersection>-183.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-183.5,-544.5,-182.5,-544.5</points>
<connection>
<GID>523</GID>
<name>IN_1</name></connection>
<intersection>-183.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-183.5,-540,-182.5,-540</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>-183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-243.5,-537,-243.5,-537</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,-509.5,-141,-509.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>-195.5 4</intersection>
<intersection>-186.5 6</intersection>
<intersection>-177.5 7</intersection>
<intersection>-168 8</intersection>
<intersection>-159 9</intersection>
<intersection>-150 10</intersection>
<intersection>-141 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-141,-510,-141,-509.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-195.5,-510,-195.5,-509.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-186.5,-510,-186.5,-509.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-177.5,-510,-177.5,-509.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-168,-510,-168,-509.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-159,-510,-159,-509.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-150,-510,-150,-509.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>-509.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-194,-543.5,-188,-543.5</points>
<connection>
<GID>511</GID>
<name>OUT</name></connection>
<connection>
<GID>524</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-199.5,-510,-199.5,-508</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-210,-508,-145,-508</points>
<intersection>-210 2</intersection>
<intersection>-199.5 0</intersection>
<intersection>-190.5 5</intersection>
<intersection>-181.5 6</intersection>
<intersection>-172 7</intersection>
<intersection>-163 8</intersection>
<intersection>-154 9</intersection>
<intersection>-145 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-210,-515.5,-210,-508</points>
<connection>
<GID>552</GID>
<name>OUT</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-145,-510,-145,-508</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-190.5,-510,-190.5,-508</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-181.5,-510,-181.5,-508</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-172,-510,-172,-508</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-163,-510,-163,-508</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-154,-510,-154,-508</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-508 1</intersection></vsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-220,-508.5,-217,-508.5</points>
<connection>
<GID>550</GID>
<name>CLK</name></connection>
<connection>
<GID>467</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>4,-542,5,-542</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>555</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>7,-542,8,-542</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<connection>
<GID>557</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>538</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>86.5,-643,89,-643</points>
<connection>
<GID>592</GID>
<name>IN_1</name></connection>
<intersection>86.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>86.5,-644.5,86.5,-643</points>
<intersection>-644.5 12</intersection>
<intersection>-643 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>80.5,-644.5,86.5,-644.5</points>
<connection>
<GID>591</GID>
<name>CLK</name></connection>
<intersection>86.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-639,82.5,-639</points>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection>
<connection>
<GID>596</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-547.5,1.5,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-547.5,4.5,-547.5</points>
<intersection>1.5 0</intersection>
<intersection>4.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-536,3,-536</points>
<connection>
<GID>555</GID>
<name>IN_1</name></connection>
<intersection>1.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-550,4.5,-547.5</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>13,-542,14,-542</points>
<connection>
<GID>566</GID>
<name>IN_1</name></connection>
<connection>
<GID>564</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>16,-542,17,-542</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<connection>
<GID>565</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-547.5,10.5,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-547.5,13.5,-547.5</points>
<intersection>10.5 0</intersection>
<intersection>13.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-536,12,-536</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-550,13.5,-547.5</points>
<connection>
<GID>562</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>22,-542,23,-542</points>
<connection>
<GID>570</GID>
<name>IN_1</name></connection>
<connection>
<GID>568</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>25,-542,26,-542</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<connection>
<GID>569</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-547.5,19.5,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-547.5,22.5,-547.5</points>
<intersection>19.5 0</intersection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-536,21,-536</points>
<connection>
<GID>568</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-550,22.5,-547.5</points>
<connection>
<GID>567</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>31.5,-542,32.5,-542</points>
<connection>
<GID>574</GID>
<name>IN_1</name></connection>
<connection>
<GID>572</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>34.5,-542,35.5,-542</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-547.5,29,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-547.5,32,-547.5</points>
<intersection>29 0</intersection>
<intersection>32 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-536,30.5,-536</points>
<connection>
<GID>572</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-550,32,-547.5</points>
<connection>
<GID>571</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>40.5,-542,41.5,-542</points>
<connection>
<GID>578</GID>
<name>IN_1</name></connection>
<connection>
<GID>576</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>43.5,-542,44.5,-542</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<connection>
<GID>577</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-547.5,38,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-547.5,41,-547.5</points>
<intersection>38 0</intersection>
<intersection>41 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-536,39.5,-536</points>
<connection>
<GID>576</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-550,41,-547.5</points>
<connection>
<GID>575</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>49.5,-542,50.5,-542</points>
<connection>
<GID>582</GID>
<name>IN_1</name></connection>
<connection>
<GID>580</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>52.5,-542,53.5,-542</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<connection>
<GID>581</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-547.5,47,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-547.5,50,-547.5</points>
<intersection>47 0</intersection>
<intersection>50 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-536,48.5,-536</points>
<connection>
<GID>580</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-550,50,-547.5</points>
<connection>
<GID>579</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58.5,-542,59.5,-542</points>
<connection>
<GID>586</GID>
<name>IN_1</name></connection>
<connection>
<GID>584</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>61.5,-542,62.5,-542</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<connection>
<GID>585</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-547.5,56,-536</points>
<intersection>-547.5 1</intersection>
<intersection>-536 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-547.5,59,-547.5</points>
<intersection>56 0</intersection>
<intersection>59 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-536,57.5,-536</points>
<connection>
<GID>584</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59,-550,59,-547.5</points>
<connection>
<GID>583</GID>
<name>OUT_0</name></connection>
<intersection>-547.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-641,89,-640</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>-640 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-640,89,-640</points>
<connection>
<GID>596</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-641,82.5,-641</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>75 14</intersection>
<intersection>81 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>81,-646.5,81,-641</points>
<intersection>-646.5 16</intersection>
<intersection>-641 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>75,-641,75,-635.5</points>
<connection>
<GID>588</GID>
<name>OUT_0</name></connection>
<intersection>-641 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>81,-646.5,87.5,-646.5</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>81 9</intersection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-550,6,-548</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-550,7.5,-550</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-550,24,-548</points>
<connection>
<GID>570</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-550,26,-550</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-550,15,-548</points>
<connection>
<GID>566</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-550,16.5,-550</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-550,33.5,-548</points>
<connection>
<GID>574</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-550,35,-550</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-550,42.5,-548</points>
<connection>
<GID>578</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-550,44,-550</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-550,51.5,-548</points>
<connection>
<GID>582</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-550,53,-550</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-550,60.5,-548</points>
<connection>
<GID>586</GID>
<name>OUT</name></connection>
<intersection>-550 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-550,62,-550</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-646.5,98.5,-642</points>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<intersection>-646.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>91.5,-646.5,98.5,-646.5</points>
<connection>
<GID>590</GID>
<name>OUT_0</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-635,97.5,-635</points>
<connection>
<GID>593</GID>
<name>clock</name></connection>
<intersection>97.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-636,97.5,-635</points>
<connection>
<GID>589</GID>
<name>OUT</name></connection>
<intersection>-635 1</intersection></vsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-216,-516.5,-216,-509.5</points>
<connection>
<GID>552</GID>
<name>IN_1</name></connection>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>-516.5 8</intersection>
<intersection>-509.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-216,-509.5,-208,-509.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-216 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-217,-516.5,-216,-516.5</points>
<connection>
<GID>698</GID>
<name>OUT_0</name></connection>
<intersection>-216 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-634,85.5,-634</points>
<connection>
<GID>593</GID>
<name>count_enable</name></connection>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-639,78.5,-623</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>-623 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-623,94.5,-623</points>
<intersection>78.5 0</intersection>
<intersection>90 3</intersection>
<intersection>94.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>94.5,-633,94.5,-623</points>
<connection>
<GID>593</GID>
<name>clear</name></connection>
<intersection>-623 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>90,-623.5,90,-623</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<intersection>-623 1</intersection></vsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-630,88.5,-629.5</points>
<connection>
<GID>593</GID>
<name>OUT_3</name></connection>
<intersection>-629.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-629.5,89,-629.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-630,91.5,-629.5</points>
<connection>
<GID>593</GID>
<name>OUT_0</name></connection>
<intersection>-629.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-629.5,91.5,-629.5</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>88.5,-619.5,97.5,-619.5</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<connection>
<GID>652</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>95,-643,102,-643</points>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<intersection>95 35</intersection>
<intersection>96.5 34</intersection>
<intersection>102 37</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>96.5,-643,96.5,-642</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<intersection>-643 6</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>95,-643,95,-642</points>
<connection>
<GID>592</GID>
<name>OUT</name></connection>
<intersection>-643 6</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>102,-643,102,-641</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>-643 6</intersection></vsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>75,-631.5,75,-631.5</points>
<connection>
<GID>563</GID>
<name>OUT_0</name></connection>
<connection>
<GID>588</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-619.5,101.5,-615.5</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<connection>
<GID>653</GID>
<name>OUT_0</name></connection>
<intersection>-615.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>101.5,-615.5,109,-615.5</points>
<intersection>101.5 0</intersection>
<intersection>109 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>109,-615.5,109,-611.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>-615.5 27</intersection></vsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>75,-627.5,75,-616.5</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<intersection>-620.5 10</intersection>
<intersection>-616.5 43</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>75,-620.5,78.5,-620.5</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>75 7</intersection>
<intersection>78.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>78.5,-620.5,78.5,-618.5</points>
<intersection>-620.5 10</intersection>
<intersection>-618.5 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>78.5,-618.5,82.5,-618.5</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>78.5 28</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>75,-616.5,79.5,-616.5</points>
<connection>
<GID>559</GID>
<name>OUT_0</name></connection>
<intersection>75 7</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-620.5,82.5,-620.5</points>
<connection>
<GID>629</GID>
<name>OUT_0</name></connection>
<connection>
<GID>652</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-612.5,79.5,-612.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<connection>
<GID>560</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>108,-633.5,214,-633.5</points>
<intersection>108 20</intersection>
<intersection>113.5 9</intersection>
<intersection>122.5 8</intersection>
<intersection>131.5 7</intersection>
<intersection>141 6</intersection>
<intersection>150 16</intersection>
<intersection>159 12</intersection>
<intersection>168 14</intersection>
<intersection>177 11</intersection>
<intersection>214 18</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>141,-633.5,141,-629.5</points>
<connection>
<GID>612</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>131.5,-633.5,131.5,-629.5</points>
<connection>
<GID>608</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>122.5,-633.5,122.5,-629.5</points>
<connection>
<GID>604</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>113.5,-633.5,113.5,-629.5</points>
<connection>
<GID>598</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>177,-633.5,177,-629.5</points>
<connection>
<GID>628</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>159,-633.5,159,-629.5</points>
<connection>
<GID>620</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>168,-633.5,168,-629.5</points>
<connection>
<GID>624</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>150,-633.5,150,-629.5</points>
<connection>
<GID>616</GID>
<name>clock</name></connection>
<intersection>-633.5 2</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>214,-633.5,214,-626</points>
<intersection>-633.5 2</intersection>
<intersection>-626 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>214,-626,215.5,-626</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>214 18</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>108,-642,108,-633.5</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<intersection>-633.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>119,-618.5,120,-618.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<connection>
<GID>599</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>122,-618.5,123,-618.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<connection>
<GID>600</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,-610,174.5,-610</points>
<intersection>107.5 27</intersection>
<intersection>120 42</intersection>
<intersection>129 34</intersection>
<intersection>138 37</intersection>
<intersection>147.5 38</intersection>
<intersection>156.5 39</intersection>
<intersection>165.5 40</intersection>
<intersection>174.5 36</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>107.5,-618.5,107.5,-610</points>
<connection>
<GID>603</GID>
<name>OUT</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>129,-612.5,129,-610</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>174.5,-612.5,174.5,-610</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>138,-612.5,138,-610</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>147.5,-612.5,147.5,-610</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>156.5,-612.5,156.5,-610</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>165.5,-612.5,165.5,-610</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>120,-612.5,120,-610</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>-610 1</intersection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-624,116.5,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-624,119.5,-624</points>
<intersection>116.5 0</intersection>
<intersection>119.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-612.5,118,-612.5</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>116.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>119.5,-626.5,119.5,-624</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>128,-618.5,129,-618.5</points>
<connection>
<GID>607</GID>
<name>IN_1</name></connection>
<connection>
<GID>605</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>131,-618.5,132,-618.5</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<connection>
<GID>606</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-624,125.5,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-624,128.5,-624</points>
<intersection>125.5 0</intersection>
<intersection>128.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-612.5,127,-612.5</points>
<connection>
<GID>605</GID>
<name>IN_1</name></connection>
<intersection>125.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-626.5,128.5,-624</points>
<connection>
<GID>604</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>137,-618.5,138,-618.5</points>
<connection>
<GID>611</GID>
<name>IN_1</name></connection>
<connection>
<GID>609</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>140,-618.5,141,-618.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<connection>
<GID>610</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-624,134.5,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-624,137.5,-624</points>
<intersection>134.5 0</intersection>
<intersection>137.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-612.5,136,-612.5</points>
<connection>
<GID>609</GID>
<name>IN_1</name></connection>
<intersection>134.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137.5,-626.5,137.5,-624</points>
<connection>
<GID>608</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>146.5,-618.5,147.5,-618.5</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<connection>
<GID>613</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>149.5,-618.5,150.5,-618.5</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<connection>
<GID>614</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-624,144,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-624,147,-624</points>
<intersection>144 0</intersection>
<intersection>147 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144,-612.5,145.5,-612.5</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<intersection>144 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>147,-626.5,147,-624</points>
<connection>
<GID>612</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155.5,-618.5,156.5,-618.5</points>
<connection>
<GID>619</GID>
<name>IN_1</name></connection>
<connection>
<GID>617</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>158.5,-618.5,159.5,-618.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<connection>
<GID>618</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-624,153,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,-624,156,-624</points>
<intersection>153 0</intersection>
<intersection>156 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153,-612.5,154.5,-612.5</points>
<connection>
<GID>617</GID>
<name>IN_1</name></connection>
<intersection>153 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>156,-626.5,156,-624</points>
<connection>
<GID>616</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>164.5,-618.5,165.5,-618.5</points>
<connection>
<GID>621</GID>
<name>OUT</name></connection>
<connection>
<GID>623</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>167.5,-618.5,168.5,-618.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<connection>
<GID>622</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-624,162,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-624,165,-624</points>
<intersection>162 0</intersection>
<intersection>165 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162,-612.5,163.5,-612.5</points>
<connection>
<GID>621</GID>
<name>IN_1</name></connection>
<intersection>162 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>165,-626.5,165,-624</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>173.5,-618.5,174.5,-618.5</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<connection>
<GID>625</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>176.5,-618.5,177.5,-618.5</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<connection>
<GID>626</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-624,171,-612.5</points>
<intersection>-624 1</intersection>
<intersection>-612.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-624,174,-624</points>
<intersection>171 0</intersection>
<intersection>174 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-612.5,172.5,-612.5</points>
<connection>
<GID>625</GID>
<name>IN_1</name></connection>
<intersection>171 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>174,-626.5,174,-624</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<intersection>-624 1</intersection></vsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-626.5,113.5,-609</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>-609 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-609,113.5,-609</points>
<connection>
<GID>630</GID>
<name>OUT_0</name></connection>
<intersection>113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-626.5,121,-624.5</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-626.5,122.5,-626.5</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-626.5,139,-624.5</points>
<connection>
<GID>611</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-626.5,141,-626.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-626.5,130,-624.5</points>
<connection>
<GID>607</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-626.5,131.5,-626.5</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-626.5,148.5,-624.5</points>
<connection>
<GID>615</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-626.5,150,-626.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-626.5,157.5,-624.5</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-626.5,159,-626.5</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-626.5,166.5,-624.5</points>
<connection>
<GID>623</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-626.5,168,-626.5</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-626.5,175.5,-624.5</points>
<connection>
<GID>627</GID>
<name>OUT</name></connection>
<intersection>-626.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-626.5,177,-626.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-612.5,176.5,-602</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>-602 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-602,176.5,-602</points>
<connection>
<GID>630</GID>
<name>OUT_7</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-612.5,167.5,-603</points>
<connection>
<GID>622</GID>
<name>IN_1</name></connection>
<intersection>-603 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-603,167.5,-603</points>
<connection>
<GID>630</GID>
<name>OUT_6</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-612.5,158.5,-604</points>
<connection>
<GID>618</GID>
<name>IN_1</name></connection>
<intersection>-604 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-604,158.5,-604</points>
<connection>
<GID>630</GID>
<name>OUT_5</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-612.5,149.5,-605</points>
<connection>
<GID>614</GID>
<name>IN_1</name></connection>
<intersection>-605 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-605,149.5,-605</points>
<connection>
<GID>630</GID>
<name>OUT_4</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-612.5,140,-606</points>
<connection>
<GID>610</GID>
<name>IN_1</name></connection>
<intersection>-606 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-606,140,-606</points>
<connection>
<GID>630</GID>
<name>OUT_3</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-612.5,131,-607</points>
<connection>
<GID>606</GID>
<name>IN_1</name></connection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-607,131,-607</points>
<connection>
<GID>630</GID>
<name>OUT_2</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>102.5,-611,102.5,-611</points>
<connection>
<GID>630</GID>
<name>clock</name></connection>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-612.5,98.5,-609</points>
<intersection>-612.5 2</intersection>
<intersection>-609 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-609,99.5,-609</points>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-612.5,98.5,-612.5</points>
<connection>
<GID>640</GID>
<name>OUT_0</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-610.5,97,-608</points>
<intersection>-610.5 1</intersection>
<intersection>-608 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-610.5,97,-610.5</points>
<connection>
<GID>639</GID>
<name>OUT_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-608,99.5,-608</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-608.5,96.5,-607</points>
<intersection>-608.5 2</intersection>
<intersection>-607 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-607,99.5,-607</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-608.5,96.5,-608.5</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-606.5,95.5,-606</points>
<intersection>-606.5 1</intersection>
<intersection>-606 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-606.5,95.5,-606.5</points>
<connection>
<GID>637</GID>
<name>OUT_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-606,99.5,-606</points>
<connection>
<GID>630</GID>
<name>IN_3</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-605,95.5,-604.5</points>
<intersection>-605 1</intersection>
<intersection>-604.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-605,99.5,-605</points>
<connection>
<GID>630</GID>
<name>IN_4</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-604.5,95.5,-604.5</points>
<connection>
<GID>636</GID>
<name>OUT_0</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-603,97.5,-600.5</points>
<intersection>-603 1</intersection>
<intersection>-600.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-603,99.5,-603</points>
<connection>
<GID>630</GID>
<name>IN_6</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-600.5,97.5,-600.5</points>
<connection>
<GID>634</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-604,96.5,-602.5</points>
<intersection>-604 2</intersection>
<intersection>-602.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-602.5,96.5,-602.5</points>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-604,99.5,-604</points>
<connection>
<GID>630</GID>
<name>IN_5</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-602,98.5,-598.5</points>
<intersection>-602 2</intersection>
<intersection>-598.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-598.5,98.5,-598.5</points>
<connection>
<GID>633</GID>
<name>OUT_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-602,99.5,-602</points>
<connection>
<GID>630</GID>
<name>IN_7</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>102.5,-600,102.5,-600</points>
<connection>
<GID>630</GID>
<name>load</name></connection>
<connection>
<GID>632</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-606,222,-602.5</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>-606 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-606,222,-606</points>
<intersection>210.5 2</intersection>
<intersection>222 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>210.5,-606,210.5,-581</points>
<connection>
<GID>515</GID>
<name>OUT</name></connection>
<intersection>-606 1</intersection></vsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-596.5,222,-594</points>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>-595.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-595.5,245,-595.5</points>
<intersection>222 0</intersection>
<intersection>245 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>245,-595.5,245,-576.5</points>
<intersection>-595.5 1</intersection>
<intersection>-576.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>245,-576.5,247,-576.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>245 2</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-588,222,-585.5</points>
<connection>
<GID>643</GID>
<name>OUT_0</name></connection>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>-587 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-587,244,-587</points>
<intersection>222 0</intersection>
<intersection>244 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>244,-587,244,-575.5</points>
<intersection>-587 3</intersection>
<intersection>-575.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>244,-575.5,247,-575.5</points>
<connection>
<GID>641</GID>
<name>IN_1</name></connection>
<intersection>244 4</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-579.5,222,-577.5</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>-578.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>222,-578.5,243,-578.5</points>
<intersection>222 0</intersection>
<intersection>243 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>243,-578.5,243,-574.5</points>
<intersection>-578.5 6</intersection>
<intersection>-574.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>243,-574.5,247,-574.5</points>
<connection>
<GID>641</GID>
<name>IN_2</name></connection>
<intersection>243 7</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-571.5,222,-570</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>-570.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-570.5,242,-570.5</points>
<intersection>222 0</intersection>
<intersection>242 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>242,-573.5,242,-570.5</points>
<intersection>-573.5 5</intersection>
<intersection>-570.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>242,-573.5,247,-573.5</points>
<connection>
<GID>641</GID>
<name>IN_3</name></connection>
<intersection>242 4</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-572.5,243,-563.5</points>
<intersection>-572.5 5</intersection>
<intersection>-563.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>243,-572.5,247,-572.5</points>
<connection>
<GID>641</GID>
<name>IN_4</name></connection>
<intersection>243 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>222,-563.5,243,-563.5</points>
<intersection>222 8</intersection>
<intersection>243 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>222,-564,222,-562.5</points>
<connection>
<GID>646</GID>
<name>OUT_0</name></connection>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-563.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-556.5,222,-555</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-555.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-555.5,244,-555.5</points>
<intersection>222 0</intersection>
<intersection>244 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>244,-571.5,244,-555.5</points>
<intersection>-571.5 5</intersection>
<intersection>-555.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>244,-571.5,247,-571.5</points>
<connection>
<GID>641</GID>
<name>IN_5</name></connection>
<intersection>244 4</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-549,222,-547.5</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-548 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>222,-548,245,-548</points>
<intersection>222 0</intersection>
<intersection>245 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>245,-570.5,245,-548</points>
<intersection>-570.5 5</intersection>
<intersection>-548 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>245,-570.5,247,-570.5</points>
<connection>
<GID>641</GID>
<name>IN_6</name></connection>
<intersection>245 4</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-541.5,222,-539</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<intersection>-539 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-539,247,-539</points>
<intersection>222 0</intersection>
<intersection>247 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>247,-569.5,247,-539</points>
<connection>
<GID>641</GID>
<name>IN_7</name></connection>
<intersection>-539 1</intersection></vsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>250,-567.5,250,-567.5</points>
<connection>
<GID>641</GID>
<name>load</name></connection>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-626.5,194.5,-582</points>
<intersection>-626.5 2</intersection>
<intersection>-582 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-582,206.5,-582</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183,-626.5,194.5,-626.5</points>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-612.5,124,-611.5</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-611.5,178.5,-611.5</points>
<connection>
<GID>655</GID>
<name>OUT_0</name></connection>
<intersection>124 0</intersection>
<intersection>133 5</intersection>
<intersection>142 6</intersection>
<intersection>151.5 7</intersection>
<intersection>160.5 8</intersection>
<intersection>169.5 9</intersection>
<intersection>178.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>178.5,-612.5,178.5,-611.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>133,-612.5,133,-611.5</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>142,-612.5,142,-611.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>151.5,-612.5,151.5,-611.5</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>160.5,-612.5,160.5,-611.5</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>169.5,-612.5,169.5,-611.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>-611.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-608.5,83.5,-608.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-595.5,63,-584.5</points>
<connection>
<GID>547</GID>
<name>IN_1</name></connection>
<intersection>-584.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19,-584.5,63,-584.5</points>
<intersection>-19 2</intersection>
<intersection>63 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-19,-608,-19,-584.5</points>
<intersection>-608 3</intersection>
<intersection>-584.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-30,-608,-19,-608</points>
<connection>
<GID>486</GID>
<name>OUT_7</name></connection>
<intersection>-19 2</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-550,-13,-532</points>
<intersection>-550 1</intersection>
<intersection>-532 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-550,-1.5,-550</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32,-532,-13,-532</points>
<connection>
<GID>475</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-536,7,-531</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<intersection>-531 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-531,7,-531</points>
<connection>
<GID>475</GID>
<name>OUT_1</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-536,16,-530</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>-530 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-530,16,-530</points>
<connection>
<GID>475</GID>
<name>OUT_2</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-536,25,-529</points>
<connection>
<GID>569</GID>
<name>IN_1</name></connection>
<intersection>-529 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-529,25,-529</points>
<connection>
<GID>475</GID>
<name>OUT_3</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-536,34.5,-528</points>
<connection>
<GID>573</GID>
<name>IN_1</name></connection>
<intersection>-528 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-528,34.5,-528</points>
<connection>
<GID>475</GID>
<name>OUT_4</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-5,-594,-5,-494</points>
<intersection>-594 59</intersection>
<intersection>-534 37</intersection>
<intersection>-494 35</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>-132,-543.5,-132,-494</points>
<intersection>-543.5 88</intersection>
<intersection>-494 35</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>-132,-494,-5,-494</points>
<intersection>-132 22</intersection>
<intersection>-5 2</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-5,-534,59.5,-534</points>
<intersection>-5 2</intersection>
<intersection>5 80</intersection>
<intersection>14 52</intersection>
<intersection>23 53</intersection>
<intersection>32.5 54</intersection>
<intersection>41.5 55</intersection>
<intersection>50.5 56</intersection>
<intersection>59.5 51</intersection></hsegment>
<vsegment>
<ID>51</ID>
<points>59.5,-536,59.5,-534</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>14,-536,14,-534</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>23,-536,23,-534</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>32.5,-536,32.5,-534</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>41.5,-536,41.5,-534</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>50.5,-536,50.5,-534</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<hsegment>
<ID>59</ID>
<points>-5,-594,61,-594</points>
<intersection>-5 2</intersection>
<intersection>6.5 60</intersection>
<intersection>15.5 74</intersection>
<intersection>24.5 75</intersection>
<intersection>34 76</intersection>
<intersection>43 77</intersection>
<intersection>52 78</intersection>
<intersection>61 73</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>6.5,-595.5,6.5,-594</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>61,-595.5,61,-594</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>15.5,-595.5,15.5,-594</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>24.5,-595.5,24.5,-594</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>34,-595.5,34,-594</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>43,-595.5,43,-594</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>52,-595.5,52,-594</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>-594 59</intersection></vsegment>
<vsegment>
<ID>80</ID>
<points>5,-536,5,-534</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<intersection>-534 37</intersection></vsegment>
<hsegment>
<ID>88</ID>
<points>-176.5,-543.5,-132,-543.5</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<intersection>-132 22</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-536,52.5,-526</points>
<connection>
<GID>581</GID>
<name>IN_1</name></connection>
<intersection>-526 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-526,52.5,-526</points>
<connection>
<GID>475</GID>
<name>OUT_6</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-536,61.5,-525</points>
<connection>
<GID>585</GID>
<name>IN_1</name></connection>
<intersection>-525 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-525,61.5,-525</points>
<connection>
<GID>475</GID>
<name>OUT_7</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-615,-12,-609.5</points>
<intersection>-615 1</intersection>
<intersection>-609.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-615,-12,-615</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12,-609.5,0,-609.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-595.5,8.5,-590.5</points>
<connection>
<GID>521</GID>
<name>IN_1</name></connection>
<intersection>-590.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-590.5,8.5,-590.5</points>
<intersection>-13 2</intersection>
<intersection>8.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-13,-614,-13,-590.5</points>
<intersection>-614 5</intersection>
<intersection>-590.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-30,-614,-13,-614</points>
<connection>
<GID>486</GID>
<name>OUT_1</name></connection>
<intersection>-13 2</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-595.5,17.5,-589.5</points>
<connection>
<GID>527</GID>
<name>IN_1</name></connection>
<intersection>-589.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-589.5,17.5,-589.5</points>
<intersection>-14 2</intersection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-14,-613,-14,-589.5</points>
<intersection>-613 3</intersection>
<intersection>-589.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-30,-613,-14,-613</points>
<connection>
<GID>486</GID>
<name>OUT_2</name></connection>
<intersection>-14 2</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-595.5,26.5,-588.5</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<intersection>-588.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-588.5,26.5,-588.5</points>
<intersection>-15 2</intersection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-15,-612,-15,-588.5</points>
<intersection>-612 3</intersection>
<intersection>-588.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-30,-612,-15,-612</points>
<connection>
<GID>486</GID>
<name>OUT_3</name></connection>
<intersection>-15 2</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-595.5,36,-587.5</points>
<connection>
<GID>535</GID>
<name>IN_1</name></connection>
<intersection>-587.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-587.5,36,-587.5</points>
<intersection>-16 2</intersection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-16,-611,-16,-587.5</points>
<intersection>-611 3</intersection>
<intersection>-587.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-30,-611,-16,-611</points>
<connection>
<GID>486</GID>
<name>OUT_4</name></connection>
<intersection>-16 2</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-595.5,45,-586.5</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>-586.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-586.5,45,-586.5</points>
<intersection>-17 2</intersection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-17,-610,-17,-586.5</points>
<intersection>-610 5</intersection>
<intersection>-586.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-30,-610,-17,-610</points>
<connection>
<GID>486</GID>
<name>OUT_5</name></connection>
<intersection>-17 2</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-595.5,54,-585.5</points>
<connection>
<GID>543</GID>
<name>IN_1</name></connection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18,-585.5,54,-585.5</points>
<intersection>-18 2</intersection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-18,-609,-18,-585.5</points>
<intersection>-609 3</intersection>
<intersection>-585.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-30,-609,-18,-609</points>
<connection>
<GID>486</GID>
<name>OUT_6</name></connection>
<intersection>-18 2</intersection></hsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-625,231.5,-547.5</points>
<intersection>-625 1</intersection>
<intersection>-602.5 4</intersection>
<intersection>-594 3</intersection>
<intersection>-585.5 10</intersection>
<intersection>-577.5 9</intersection>
<intersection>-570 8</intersection>
<intersection>-562.5 11</intersection>
<intersection>-555 12</intersection>
<intersection>-547.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221.5,-625,250,-625</points>
<connection>
<GID>667</GID>
<name>OUT</name></connection>
<intersection>231.5 0</intersection>
<intersection>250 14</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>225,-594,231.5,-594</points>
<connection>
<GID>643</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>225,-602.5,231.5,-602.5</points>
<connection>
<GID>642</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>225,-547.5,231.5,-547.5</points>
<connection>
<GID>649</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>225,-570,231.5,-570</points>
<connection>
<GID>646</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>225,-577.5,231.5,-577.5</points>
<connection>
<GID>645</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>225,-585.5,231.5,-585.5</points>
<connection>
<GID>644</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>225,-562.5,231.5,-562.5</points>
<connection>
<GID>647</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>225,-555,231.5,-555</points>
<connection>
<GID>648</GID>
<name>clock</name></connection>
<intersection>231.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>250,-625,250,-582.5</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-625 1</intersection></vsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-612.5,122,-608</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>-608 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-608,122,-608</points>
<connection>
<GID>630</GID>
<name>OUT_1</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-578.5,250,-578.5</points>
<connection>
<GID>641</GID>
<name>clock</name></connection>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-192,-354.5,-192,-354.5</points>
<connection>
<GID>669</GID>
<name>N_in0</name></connection>
<connection>
<GID>794</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-192,-358.5,-192,-358.5</points>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection>
<connection>
<GID>670</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>-243.5,-533,-243.5,-525.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>807</GID>
<name>OUT_0</name></connection>
<intersection>-526 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-243.5,-526,-240,-526</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>-243.5 7</intersection>
<intersection>-240 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-240,-526,-240,-524</points>
<intersection>-526 10</intersection>
<intersection>-524 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>-240,-524,-236,-524</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>-240 28</intersection></hsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-192,-381.5,-192,-381.5</points>
<connection>
<GID>741</GID>
<name>OUT</name></connection>
<connection>
<GID>671</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-236,-526,-236,-526</points>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 1>
<page 2>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 2>
<page 3>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 3>
<page 4>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 4>
<page 5>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 5>
<page 6>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 6>
<page 7>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 7>
<page 8>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 8>
<page 9>
<PageViewport>-10.6032,1477.97,1383.4,775.97</PageViewport></page 9></circuit>