<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 0>
<page 1>
<PageViewport>-12.6454,-182.891,161.605,-270.641</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>77,151.5</position>
<gparam>LABEL_TEXT Bidirectional Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>88.5,60</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>91,88.5</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>230.5,-291.5</position>
<input>
<ID>N_in0</ID>276 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>BE_JKFF_LOW</type>
<position>82,127.5</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>12 </output>
<input>
<ID>clock</ID>3 </input>
<output>
<ID>nQ</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>27,-12</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>155.5,-502</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>27,-27.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>BE_JKFF_LOW</type>
<position>105,127.5</position>
<input>
<ID>J</ID>16 </input>
<input>
<ID>K</ID>16 </input>
<output>
<ID>Q</ID>19 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>57,-20</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>148.5,-501.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>57,-26.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>67,127.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>46.5,-20</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>230.5,-303.5</position>
<input>
<ID>N_in0</ID>279 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>46,-26.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>59,128</position>
<gparam>LABEL_TEXT Up/Down</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>38,-19</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>230.5,-295.5</position>
<input>
<ID>N_in0</ID>277 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>75,137.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>230.5,-299.5</position>
<input>
<ID>N_in0</ID>278 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>69,138</position>
<gparam>LABEL_TEXT Logic1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>230.5,-307.5</position>
<input>
<ID>N_in0</ID>280 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>67.5,117.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>230.5,-311.5</position>
<input>
<ID>N_in0</ID>281 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>61,118</position>
<gparam>LABEL_TEXT Toggle</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>230.5,-315.5</position>
<input>
<ID>N_in0</ID>282 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>102,-16</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>102.5,-31.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>125.5,-24</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>89,133.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>121.5,-24</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>230.5,-319.5</position>
<input>
<ID>N_in0</ID>283 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-23</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>88,121</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>28.5,-7</position>
<gparam>LABEL_TEXT 1:2 Demux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>102.5,-33.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>102.5,-35.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>102.5,-37.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>102.5,-39.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>102.5,-41.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>102.5,-43.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>102.5,-45.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>236,-230</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AE_SMALL_INVERTER</type>
<position>82.5,120</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>121.5,-28</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>121.5,-32</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>121.5,-36</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>121.5,-40</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>121.5,-44</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>236.5,-266</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>121.5,-48</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>121.5,-52</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR2</type>
<position>95,129.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>236,-304.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>85,140.5</position>
<input>
<ID>N_in2</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AE_OR2</type>
<position>226,-251.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>108,139.5</position>
<input>
<ID>N_in2</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AE_OR2</type>
<position>226,-255.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>269 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>125.5,-36</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>125.5,-28</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>125.5,-32</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>125.5,-40</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>125.5,-44</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>125.5,-48</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>125.5,-52</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>125.5,-58</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>121.5,-58</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>121.5,-62</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>121.5,-66</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>121.5,-70</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>121.5,-74</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>121.5,-78</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>121.5,-82</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>121.5,-86</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>125.5,-70</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>125.5,-62</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>125.5,-66</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>125.5,-74</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>125.5,-78</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>125.5,-82</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>125.5,-86</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-27</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-31</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-35</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-39</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-43</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-47</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_SMALL_INVERTER</type>
<position>116.5,-51</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>104.5,-8.5</position>
<gparam>LABEL_TEXT 1:2 Demux with 8bit input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>84.5,144.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>88,-37</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>183,-14</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>108,143.5</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>215.5,-22</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND2</type>
<position>211.5,-22</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-21</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>226,-259.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>270 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_OR2</type>
<position>226,-263.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>BE_JKFF_LOW</type>
<position>234,95</position>
<input>
<ID>J</ID>27 </input>
<input>
<ID>K</ID>27 </input>
<output>
<ID>Q</ID>39 </output>
<input>
<ID>clock</ID>28 </input>
<output>
<ID>nQ</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>BE_JKFF_LOW</type>
<position>257,95</position>
<input>
<ID>J</ID>123 </input>
<input>
<ID>K</ID>123 </input>
<output>
<ID>Q</ID>124 </output>
<input>
<ID>clock</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_OR2</type>
<position>226,-267.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_OR2</type>
<position>226,-271.5</position>
<input>
<ID>IN_0</ID>265 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>227,105</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>211.5,-26</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND2</type>
<position>211.5,-30</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>211.5,-34</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>211.5,-38</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>211.5,-42</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>211.5,-46</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>211.5,-50</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>215.5,-34</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>215.5,-26</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>215.5,-30</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>215.5,-38</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>215.5,-42</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>GA_LED</type>
<position>215.5,-46</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>215.5,-50</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>215.5,-56</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>211.5,-56</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>211.5,-60</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_AND2</type>
<position>211.5,-64</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND2</type>
<position>211.5,-68</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>211.5,-72</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>211.5,-76</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND2</type>
<position>211.5,-80</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>211.5,-84</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>215.5,-68</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>215.5,-60</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>GA_LED</type>
<position>215.5,-64</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>215.5,-72</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>GA_LED</type>
<position>215.5,-76</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>GA_LED</type>
<position>215.5,-80</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>215.5,-84</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-25</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-29</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-33</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-37</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-41</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-45</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-49</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>194.5,-6.5</position>
<gparam>LABEL_TEXT 2 8bit 1:2 Demux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>177.5,-35</position>
<gparam>LABEL_TEXT ~C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_TOGGLE</type>
<position>192.5,-99</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>145</ID>
<type>GA_LED</type>
<position>215.5,-91.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND2</type>
<position>211.5,-91.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-90.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>192.5,-101</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>192.5,-103</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>192.5,-105</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>192.5,-107</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>192.5,-109</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>192.5,-111</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>192.5,-113</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>211.5,-95.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>211.5,-99.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>211.5,-103.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_AND2</type>
<position>211.5,-107.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>211.5,-111.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND2</type>
<position>211.5,-115.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>211.5,-119.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>215.5,-103.5</position>
<input>
<ID>N_in0</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>215.5,-95.5</position>
<input>
<ID>N_in0</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>GA_LED</type>
<position>215.5,-99.5</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>215.5,-107.5</position>
<input>
<ID>N_in0</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>215.5,-111.5</position>
<input>
<ID>N_in0</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>215.5,-115.5</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>GA_LED</type>
<position>215.5,-119.5</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>215.5,-125.5</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>211.5,-125.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND2</type>
<position>211.5,-129.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND2</type>
<position>211.5,-133.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>211.5,-137.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>211.5,-141.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>211.5,-145.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>211.5,-149.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>211.5,-153.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>215.5,-137.5</position>
<input>
<ID>N_in0</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>GA_LED</type>
<position>215.5,-129.5</position>
<input>
<ID>N_in0</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>GA_LED</type>
<position>215.5,-133.5</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>GA_LED</type>
<position>215.5,-141.5</position>
<input>
<ID>N_in0</ID>110 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>215.5,-145.5</position>
<input>
<ID>N_in0</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>GA_LED</type>
<position>215.5,-149.5</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>215.5,-153.5</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-94.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-98.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-102.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-106.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-110.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-114.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_SMALL_INVERTER</type>
<position>206.5,-118.5</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>178,-104.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>221,105.5</position>
<gparam>LABEL_TEXT Logic1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>173,-14.5</position>
<gparam>LABEL_TEXT Flip</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AE_OR2</type>
<position>226,-275.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_OR2</type>
<position>226,-279.5</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>246 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_AND2</type>
<position>241,101</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>240,88.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_SMALL_INVERTER</type>
<position>234.5,87.5</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR2</type>
<position>247,97</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>GA_LED</type>
<position>237,108</position>
<input>
<ID>N_in2</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>GA_LED</type>
<position>260,107</position>
<input>
<ID>N_in2</ID>124 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>236.5,112</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-29.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-31.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-33.5</position>
<input>
<ID>IN_0</ID>171 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-35.5</position>
<input>
<ID>IN_0</ID>176 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-37.5</position>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>209</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-39.5</position>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-41.5</position>
<input>
<ID>IN_0</ID>174 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-43.5</position>
<input>
<ID>IN_0</ID>175 </input>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>259.5,111</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>207.5,80.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>139.5,-196</position>
<gparam>LABEL_TEXT Flip</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_TOGGLE</type>
<position>186,79</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>186,75</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>173,87.5</position>
<gparam>LABEL_TEXT Thermometer signals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>178.5,79.5</position>
<gparam>LABEL_TEXT Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>177.5,75.5</position>
<gparam>LABEL_TEXT Increase/Decrease</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>196,116</position>
<gparam>LABEL_TEXT Counter and register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AE_SMALL_INVERTER</type>
<position>218.5,87.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>208,90</position>
<gparam>LABEL_TEXT Load/Count</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_TOGGLE</type>
<position>144.5,-197.5</position>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>224</ID>
<type>GA_LED</type>
<position>202,-204.5</position>
<input>
<ID>N_in0</ID>134 </input>
<input>
<ID>N_in1</ID>252 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_TOGGLE</type>
<position>213.5,89.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>226</ID>
<type>AE_REGISTER8</type>
<position>218.5,79.5</position>
<output>
<ID>carry_out</ID>28 </output>
<input>
<ID>clock</ID>125 </input>
<input>
<ID>count_enable</ID>128 </input>
<input>
<ID>count_up</ID>129 </input>
<input>
<ID>load</ID>126 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 144</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>198,-204.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-203.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>198,-208.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>198,-212.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>BE_JKFF_LOW</type>
<position>176.5,-468.5</position>
<input>
<ID>J</ID>130 </input>
<input>
<ID>K</ID>130 </input>
<output>
<ID>Q</ID>1193 </output>
<input>
<ID>clear</ID>1 </input>
<input>
<ID>clock</ID>131 </input>
<output>
<ID>nQ</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>232</ID>
<type>BE_JKFF_LOW</type>
<position>199.5,-468.5</position>
<input>
<ID>J</ID>137 </input>
<input>
<ID>K</ID>137 </input>
<output>
<ID>Q</ID>1119 </output>
<input>
<ID>clear</ID>1 </input>
<input>
<ID>clock</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>169.5,-458.5</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>163,-458</position>
<gparam>LABEL_TEXT Logic1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_AND2</type>
<position>183.5,-462.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>1193 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>182.5,-475</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_SMALL_INVERTER</type>
<position>177,-476</position>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_OR2</type>
<position>189.5,-466.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>198,-216.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>198,-220.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>181,-417.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>198,-224.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>150,-483</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_TOGGLE</type>
<position>128.5,-484.5</position>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_TOGGLE</type>
<position>128.5,-488.5</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>115.5,-476</position>
<gparam>LABEL_TEXT Thermometer signals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>124,-484</position>
<gparam>LABEL_TEXT Update</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>120,-488</position>
<gparam>LABEL_TEXT Increase/Decrease</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_AND2</type>
<position>198,-228.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AE_SMALL_INVERTER</type>
<position>161,-476</position>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>141 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>152,-474</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>156,-474</position>
<output>
<ID>OUT_0</ID>140 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_REGISTER8</type>
<position>161,-484</position>
<output>
<ID>OUT_0</ID>150 </output>
<output>
<ID>OUT_1</ID>149 </output>
<output>
<ID>OUT_2</ID>148 </output>
<output>
<ID>OUT_3</ID>147 </output>
<output>
<ID>OUT_4</ID>146 </output>
<output>
<ID>OUT_5</ID>145 </output>
<output>
<ID>OUT_6</ID>144 </output>
<output>
<ID>OUT_7</ID>143 </output>
<output>
<ID>carry_out</ID>131 </output>
<input>
<ID>clear</ID>1 </input>
<input>
<ID>clock</ID>139 </input>
<input>
<ID>count_enable</ID>141 </input>
<input>
<ID>count_up</ID>142 </input>
<input>
<ID>load</ID>140 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>198,-232.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>GA_LED</type>
<position>202,-216.5</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>255 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>202,-414</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>GA_LED</type>
<position>202,-208.5</position>
<input>
<ID>N_in0</ID>190 </input>
<input>
<ID>N_in1</ID>253 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>GA_LED</type>
<position>202,-212.5</position>
<input>
<ID>N_in0</ID>189 </input>
<input>
<ID>N_in1</ID>254 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>GA_LED</type>
<position>202,-220.5</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>256 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>GA_LED</type>
<position>202,-224.5</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>257 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>202,-228.5</position>
<input>
<ID>N_in0</ID>194 </input>
<input>
<ID>N_in1</ID>258 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_TOGGLE</type>
<position>189,-29.5</position>
<output>
<ID>OUT_0</ID>169 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_TOGGLE</type>
<position>189,-31.5</position>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_TOGGLE</type>
<position>189,-33.5</position>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>189,-35.5</position>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_TOGGLE</type>
<position>189,-38</position>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_TOGGLE</type>
<position>189,-39.5</position>
<output>
<ID>OUT_0</ID>173 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_TOGGLE</type>
<position>189,-41.5</position>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_TOGGLE</type>
<position>189,-43.5</position>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>270</ID>
<type>GA_LED</type>
<position>202,-232.5</position>
<input>
<ID>N_in0</ID>195 </input>
<input>
<ID>N_in1</ID>259 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>GA_LED</type>
<position>202,-238.5</position>
<input>
<ID>N_in0</ID>196 </input>
<input>
<ID>N_in1</ID>260 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AA_AND2</type>
<position>198,-238.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_AND2</type>
<position>198,-242.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_AND2</type>
<position>198,-246.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>AA_AND2</type>
<position>198,-250.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>198,-254.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>198,-258.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>198,-262.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>198,-266.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>GA_LED</type>
<position>202,-250.5</position>
<input>
<ID>N_in0</ID>199 </input>
<input>
<ID>N_in1</ID>263 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>202,-242.5</position>
<input>
<ID>N_in0</ID>198 </input>
<input>
<ID>N_in1</ID>261 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>GA_LED</type>
<position>202,-246.5</position>
<input>
<ID>N_in0</ID>197 </input>
<input>
<ID>N_in1</ID>262 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>GA_LED</type>
<position>202,-254.5</position>
<input>
<ID>N_in0</ID>200 </input>
<input>
<ID>N_in1</ID>264 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>GA_LED</type>
<position>202,-258.5</position>
<input>
<ID>N_in0</ID>201 </input>
<input>
<ID>N_in1</ID>265 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>GA_LED</type>
<position>202,-262.5</position>
<input>
<ID>N_in0</ID>202 </input>
<input>
<ID>N_in1</ID>266 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>GA_LED</type>
<position>202,-266.5</position>
<input>
<ID>N_in0</ID>203 </input>
<input>
<ID>N_in1</ID>267 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-207.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-211.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-215.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-219.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-223.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>292</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-227.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>293</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-231.5</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>168,-184.5</position>
<gparam>LABEL_TEXT RGB Selector</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>GA_LED</type>
<position>202,-274</position>
<input>
<ID>N_in0</ID>213 </input>
<input>
<ID>N_in1</ID>268 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>198,-274</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-273</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND2</type>
<position>198,-278</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>198,-282</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>198,-286</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND2</type>
<position>198,-290</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>198,-294</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_AND2</type>
<position>198,-298</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>198,-302</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>GA_LED</type>
<position>202,-286</position>
<input>
<ID>N_in0</ID>223 </input>
<input>
<ID>N_in1</ID>271 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>GA_LED</type>
<position>202,-278</position>
<input>
<ID>N_in0</ID>222 </input>
<input>
<ID>N_in1</ID>269 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>GA_LED</type>
<position>202,-282</position>
<input>
<ID>N_in0</ID>221 </input>
<input>
<ID>N_in1</ID>270 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>GA_LED</type>
<position>202,-290</position>
<input>
<ID>N_in0</ID>224 </input>
<input>
<ID>N_in1</ID>272 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>GA_LED</type>
<position>202,-294</position>
<input>
<ID>N_in0</ID>225 </input>
<input>
<ID>N_in1</ID>273 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>GA_LED</type>
<position>202,-298</position>
<input>
<ID>N_in0</ID>226 </input>
<input>
<ID>N_in1</ID>274 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>GA_LED</type>
<position>202,-302</position>
<input>
<ID>N_in0</ID>227 </input>
<input>
<ID>N_in1</ID>275 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>GA_LED</type>
<position>202,-308</position>
<input>
<ID>N_in0</ID>228 </input>
<input>
<ID>N_in1</ID>276 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>198,-308</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>212 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AA_AND2</type>
<position>198,-312</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_AND2</type>
<position>198,-316</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>198,-320</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_AND2</type>
<position>198,-324</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_AND2</type>
<position>198,-328</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>198,-332</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>198,-336</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>GA_LED</type>
<position>202,-320</position>
<input>
<ID>N_in0</ID>231 </input>
<input>
<ID>N_in1</ID>279 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>GA_LED</type>
<position>202,-312</position>
<input>
<ID>N_in0</ID>230 </input>
<input>
<ID>N_in1</ID>277 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>GA_LED</type>
<position>202,-316</position>
<input>
<ID>N_in0</ID>229 </input>
<input>
<ID>N_in1</ID>278 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>AA_TOGGLE</type>
<position>67,58.5</position>
<output>
<ID>OUT_0</ID>312 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>325</ID>
<type>GA_LED</type>
<position>202,-324</position>
<input>
<ID>N_in0</ID>232 </input>
<input>
<ID>N_in1</ID>280 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_TOGGLE</type>
<position>67,54.5</position>
<output>
<ID>OUT_0</ID>1212 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>327</ID>
<type>GA_LED</type>
<position>202,-328</position>
<input>
<ID>N_in0</ID>233 </input>
<input>
<ID>N_in1</ID>281 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>AA_LABEL</type>
<position>54,67</position>
<gparam>LABEL_TEXT Thermometer signals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>GA_LED</type>
<position>202,-332</position>
<input>
<ID>N_in0</ID>234 </input>
<input>
<ID>N_in1</ID>282 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>330</ID>
<type>AA_LABEL</type>
<position>59.5,59</position>
<gparam>LABEL_TEXT Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>331</ID>
<type>AA_LABEL</type>
<position>58.5,55</position>
<gparam>LABEL_TEXT Increase/Decrease</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>GA_LED</type>
<position>202,-336</position>
<input>
<ID>N_in0</ID>235 </input>
<input>
<ID>N_in1</ID>283 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>333</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-277</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-281</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-285</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-289</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-293</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-297</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_SMALL_INVERTER</type>
<position>193,-301</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>340</ID>
<type>GA_LED</type>
<position>230,-215</position>
<input>
<ID>N_in0</ID>252 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>341</ID>
<type>GA_LED</type>
<position>230,-227</position>
<input>
<ID>N_in0</ID>255 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>GA_LED</type>
<position>230,-219</position>
<input>
<ID>N_in0</ID>253 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>GA_LED</type>
<position>230,-223</position>
<input>
<ID>N_in0</ID>254 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>344</ID>
<type>GA_LED</type>
<position>230,-231</position>
<input>
<ID>N_in0</ID>256 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>345</ID>
<type>GA_LED</type>
<position>230,-235</position>
<input>
<ID>N_in0</ID>257 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>GA_LED</type>
<position>230,-239</position>
<input>
<ID>N_in0</ID>258 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>GA_LED</type>
<position>230,-243</position>
<input>
<ID>N_in0</ID>259 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>GA_LED</type>
<position>230,-251.5</position>
<input>
<ID>N_in0</ID>244 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>230,-263.5</position>
<input>
<ID>N_in0</ID>248 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>230,-255.5</position>
<input>
<ID>N_in0</ID>245 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>GA_LED</type>
<position>230,-259.5</position>
<input>
<ID>N_in0</ID>247 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>GA_LED</type>
<position>230,-267.5</position>
<input>
<ID>N_in0</ID>249 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>353</ID>
<type>GA_LED</type>
<position>230,-271.5</position>
<input>
<ID>N_in0</ID>250 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>GA_LED</type>
<position>230,-275.5</position>
<input>
<ID>N_in0</ID>251 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>GA_LED</type>
<position>230,-279.5</position>
<input>
<ID>N_in0</ID>246 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>152,-204.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>376</ID>
<type>DA_FROM</type>
<position>164,-206.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_LABEL</type>
<position>153.5,-216.5</position>
<gparam>LABEL_TEXT ~C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>378</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-206.5</position>
<input>
<ID>IN_0</ID>293 </input>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>379</ID>
<type>DA_FROM</type>
<position>164,-210.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-210.5</position>
<input>
<ID>IN_0</ID>294 </input>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>381</ID>
<type>DA_FROM</type>
<position>164,-214.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_LABEL</type>
<position>64.5,86.5</position>
<gparam>LABEL_TEXT Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>383</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-214.5</position>
<input>
<ID>IN_0</ID>295 </input>
<output>
<ID>OUT_0</ID>303 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>164,-218.5</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-218.5</position>
<input>
<ID>IN_0</ID>296 </input>
<output>
<ID>OUT_0</ID>304 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>164,-222.5</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>387</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-222.5</position>
<input>
<ID>IN_0</ID>297 </input>
<output>
<ID>OUT_0</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>164,-226.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>389</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-226.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>164,-230.5</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>391</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-230.5</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>392</ID>
<type>DA_FROM</type>
<position>164,-234.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>393</ID>
<type>AE_SMALL_INVERTER</type>
<position>168,-234.5</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>307 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AE_SMALL_INVERTER</type>
<position>99.5,67</position>
<input>
<ID>IN_0</ID>322 </input>
<output>
<ID>OUT_0</ID>1210 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>395</ID>
<type>AE_OR2</type>
<position>173,-205.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>301 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_LABEL</type>
<position>89,69.5</position>
<gparam>LABEL_TEXT Load/Count</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>AE_OR2</type>
<position>173,-209.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>302 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>398</ID>
<type>AE_OR2</type>
<position>173,-213.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>303 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>AE_OR2</type>
<position>173,-217.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>173,-221.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>305 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>AE_OR2</type>
<position>173,-229.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>306 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>AE_OR2</type>
<position>173,-233.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AE_SMALL_INVERTER</type>
<position>156,-204.5</position>
<input>
<ID>IN_0</ID>308 </input>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>161.5,-274</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>167.5,-276</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_LABEL</type>
<position>158,-286.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>167.5,-280</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>408</ID>
<type>DA_FROM</type>
<position>167.5,-284</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_LABEL</type>
<position>133,-424</position>
<gparam>LABEL_TEXT Complete Circuit</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>167.5,-288</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>167.5,-292</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>167.5,-296</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>167.5,-300</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>167.5,-304</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>415</ID>
<type>AE_OR2</type>
<position>172.5,-275</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>311 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>AE_OR2</type>
<position>172.5,-279</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>AE_OR2</type>
<position>172.5,-283</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AE_OR2</type>
<position>172.5,-287</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>315 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AE_OR2</type>
<position>172.5,-291</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>316 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>420</ID>
<type>AE_OR2</type>
<position>172.5,-295</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>421</ID>
<type>AE_OR2</type>
<position>172.5,-299</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>422</ID>
<type>AE_OR2</type>
<position>172.5,-303</position>
<input>
<ID>IN_0</ID>310 </input>
<input>
<ID>IN_1</ID>317 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>34.5,-249</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>644</ID>
<type>AA_LABEL</type>
<position>260,-12</position>
<gparam>LABEL_TEXT Flip</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>645</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-27</position>
<input>
<ID>IN_0</ID>611 </input>
<output>
<ID>OUT_0</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-29</position>
<input>
<ID>IN_0</ID>610 </input>
<output>
<ID>OUT_0</ID>548 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-31</position>
<input>
<ID>IN_0</ID>614 </input>
<output>
<ID>OUT_0</ID>549 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>648</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-33</position>
<input>
<ID>IN_0</ID>617 </input>
<output>
<ID>OUT_0</ID>550 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>649</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-35</position>
<input>
<ID>IN_0</ID>612 </input>
<output>
<ID>OUT_0</ID>551 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-37</position>
<input>
<ID>IN_0</ID>613 </input>
<output>
<ID>OUT_0</ID>552 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>651</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-39</position>
<input>
<ID>IN_0</ID>616 </input>
<output>
<ID>OUT_0</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>652</ID>
<type>AE_SMALL_INVERTER</type>
<position>280,-41</position>
<input>
<ID>IN_0</ID>615 </input>
<output>
<ID>OUT_0</ID>554 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>653</ID>
<type>AA_TOGGLE</type>
<position>270,-11.5</position>
<output>
<ID>OUT_0</ID>603 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>654</ID>
<type>GA_LED</type>
<position>302.5,-19.5</position>
<input>
<ID>N_in0</ID>547 </input>
<input>
<ID>N_in1</ID>626 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>655</ID>
<type>AA_AND2</type>
<position>298.5,-19.5</position>
<input>
<ID>IN_0</ID>545 </input>
<input>
<ID>IN_1</ID>546 </input>
<output>
<ID>OUT</ID>547 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-18.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>545 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_AND2</type>
<position>298.5,-23.5</position>
<input>
<ID>IN_0</ID>576 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>AA_AND2</type>
<position>298.5,-27.5</position>
<input>
<ID>IN_0</ID>575 </input>
<input>
<ID>IN_1</ID>549 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_AND2</type>
<position>298.5,-31.5</position>
<input>
<ID>IN_0</ID>574 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>660</ID>
<type>AA_AND2</type>
<position>298.5,-35.5</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>551 </input>
<output>
<ID>OUT</ID>558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>661</ID>
<type>AA_AND2</type>
<position>298.5,-39.5</position>
<input>
<ID>IN_0</ID>572 </input>
<input>
<ID>IN_1</ID>552 </input>
<output>
<ID>OUT</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_AND2</type>
<position>298.5,-43.5</position>
<input>
<ID>IN_0</ID>571 </input>
<input>
<ID>IN_1</ID>553 </input>
<output>
<ID>OUT</ID>560 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>AA_AND2</type>
<position>298.5,-47.5</position>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>554 </input>
<output>
<ID>OUT</ID>561 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>664</ID>
<type>GA_LED</type>
<position>302.5,-31.5</position>
<input>
<ID>N_in0</ID>557 </input>
<input>
<ID>N_in1</ID>629 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>665</ID>
<type>GA_LED</type>
<position>302.5,-23.5</position>
<input>
<ID>N_in0</ID>556 </input>
<input>
<ID>N_in1</ID>627 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>666</ID>
<type>GA_LED</type>
<position>302.5,-27.5</position>
<input>
<ID>N_in0</ID>555 </input>
<input>
<ID>N_in1</ID>628 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>667</ID>
<type>GA_LED</type>
<position>302.5,-35.5</position>
<input>
<ID>N_in0</ID>558 </input>
<input>
<ID>N_in1</ID>630 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>668</ID>
<type>GA_LED</type>
<position>302.5,-39.5</position>
<input>
<ID>N_in0</ID>559 </input>
<input>
<ID>N_in1</ID>631 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>669</ID>
<type>GA_LED</type>
<position>302.5,-43.5</position>
<input>
<ID>N_in0</ID>560 </input>
<input>
<ID>N_in1</ID>632 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>670</ID>
<type>GA_LED</type>
<position>302.5,-47.5</position>
<input>
<ID>N_in0</ID>561 </input>
<input>
<ID>N_in1</ID>633 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>671</ID>
<type>GA_LED</type>
<position>302.5,-53.5</position>
<input>
<ID>N_in0</ID>562 </input>
<input>
<ID>N_in1</ID>634 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>672</ID>
<type>AA_AND2</type>
<position>298.5,-53.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>546 </input>
<output>
<ID>OUT</ID>562 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>673</ID>
<type>AA_AND2</type>
<position>298.5,-57.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>564 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>674</ID>
<type>AA_AND2</type>
<position>298.5,-61.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>549 </input>
<output>
<ID>OUT</ID>563 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_AND2</type>
<position>298.5,-65.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>676</ID>
<type>AA_AND2</type>
<position>298.5,-69.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>551 </input>
<output>
<ID>OUT</ID>566 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>677</ID>
<type>AA_AND2</type>
<position>298.5,-73.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>552 </input>
<output>
<ID>OUT</ID>567 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>678</ID>
<type>AA_AND2</type>
<position>298.5,-77.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>553 </input>
<output>
<ID>OUT</ID>568 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>679</ID>
<type>AA_AND2</type>
<position>298.5,-81.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>554 </input>
<output>
<ID>OUT</ID>569 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>680</ID>
<type>GA_LED</type>
<position>302.5,-65.5</position>
<input>
<ID>N_in0</ID>565 </input>
<input>
<ID>N_in1</ID>637 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>681</ID>
<type>GA_LED</type>
<position>302.5,-57.5</position>
<input>
<ID>N_in0</ID>564 </input>
<input>
<ID>N_in1</ID>635 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>682</ID>
<type>GA_LED</type>
<position>302.5,-61.5</position>
<input>
<ID>N_in0</ID>563 </input>
<input>
<ID>N_in1</ID>636 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>683</ID>
<type>GA_LED</type>
<position>302.5,-69.5</position>
<input>
<ID>N_in0</ID>566 </input>
<input>
<ID>N_in1</ID>638 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>684</ID>
<type>GA_LED</type>
<position>302.5,-73.5</position>
<input>
<ID>N_in0</ID>567 </input>
<input>
<ID>N_in1</ID>639 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>685</ID>
<type>GA_LED</type>
<position>302.5,-77.5</position>
<input>
<ID>N_in0</ID>568 </input>
<input>
<ID>N_in1</ID>640 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>686</ID>
<type>GA_LED</type>
<position>302.5,-81.5</position>
<input>
<ID>N_in0</ID>569 </input>
<input>
<ID>N_in1</ID>641 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>687</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-22.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>576 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>688</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-26.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>575 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>689</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-30.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-34.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-38.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>572 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>692</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-42.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>693</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-46.5</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>570 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>694</ID>
<type>AA_LABEL</type>
<position>281,-3.5</position>
<gparam>LABEL_TEXT RG/GB Flipper</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>696</ID>
<type>AA_TOGGLE</type>
<position>279.5,-96.5</position>
<output>
<ID>OUT_0</ID>578 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>697</ID>
<type>GA_LED</type>
<position>302.5,-89</position>
<input>
<ID>N_in0</ID>579 </input>
<input>
<ID>N_in1</ID>642 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>698</ID>
<type>AA_AND2</type>
<position>298.5,-89</position>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>578 </input>
<output>
<ID>OUT</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>699</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-88</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>577 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>700</ID>
<type>AA_TOGGLE</type>
<position>279.5,-98.5</position>
<output>
<ID>OUT_0</ID>580 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_TOGGLE</type>
<position>279.5,-100.5</position>
<output>
<ID>OUT_0</ID>581 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>702</ID>
<type>AA_TOGGLE</type>
<position>279.5,-102.5</position>
<output>
<ID>OUT_0</ID>582 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>703</ID>
<type>AA_TOGGLE</type>
<position>279.5,-104.5</position>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>704</ID>
<type>AA_TOGGLE</type>
<position>279.5,-106.5</position>
<output>
<ID>OUT_0</ID>584 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>705</ID>
<type>AA_TOGGLE</type>
<position>279.5,-108.5</position>
<output>
<ID>OUT_0</ID>585 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>706</ID>
<type>AA_TOGGLE</type>
<position>279.5,-110.5</position>
<output>
<ID>OUT_0</ID>586 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>707</ID>
<type>AA_AND2</type>
<position>298.5,-93</position>
<input>
<ID>IN_0</ID>609 </input>
<input>
<ID>IN_1</ID>580 </input>
<output>
<ID>OUT</ID>588 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>708</ID>
<type>AA_AND2</type>
<position>298.5,-97</position>
<input>
<ID>IN_0</ID>608 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>587 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>AA_AND2</type>
<position>298.5,-101</position>
<input>
<ID>IN_0</ID>607 </input>
<input>
<ID>IN_1</ID>582 </input>
<output>
<ID>OUT</ID>589 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_AND2</type>
<position>298.5,-105</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>583 </input>
<output>
<ID>OUT</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>711</ID>
<type>AA_AND2</type>
<position>298.5,-109</position>
<input>
<ID>IN_0</ID>605 </input>
<input>
<ID>IN_1</ID>584 </input>
<output>
<ID>OUT</ID>591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>712</ID>
<type>AA_AND2</type>
<position>298.5,-113</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>592 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>713</ID>
<type>AA_AND2</type>
<position>298.5,-117</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>586 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>714</ID>
<type>GA_LED</type>
<position>302.5,-101</position>
<input>
<ID>N_in0</ID>589 </input>
<input>
<ID>N_in1</ID>645 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>715</ID>
<type>GA_LED</type>
<position>302.5,-93</position>
<input>
<ID>N_in0</ID>588 </input>
<input>
<ID>N_in1</ID>643 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>716</ID>
<type>GA_LED</type>
<position>302.5,-97</position>
<input>
<ID>N_in0</ID>587 </input>
<input>
<ID>N_in1</ID>644 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>717</ID>
<type>GA_LED</type>
<position>302.5,-105</position>
<input>
<ID>N_in0</ID>590 </input>
<input>
<ID>N_in1</ID>646 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>718</ID>
<type>GA_LED</type>
<position>302.5,-109</position>
<input>
<ID>N_in0</ID>591 </input>
<input>
<ID>N_in1</ID>647 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>719</ID>
<type>GA_LED</type>
<position>302.5,-113</position>
<input>
<ID>N_in0</ID>592 </input>
<input>
<ID>N_in1</ID>648 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>720</ID>
<type>GA_LED</type>
<position>302.5,-117</position>
<input>
<ID>N_in0</ID>593 </input>
<input>
<ID>N_in1</ID>649 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>721</ID>
<type>GA_LED</type>
<position>302.5,-123</position>
<input>
<ID>N_in0</ID>594 </input>
<input>
<ID>N_in1</ID>650 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>722</ID>
<type>AA_AND2</type>
<position>298.5,-123</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>578 </input>
<output>
<ID>OUT</ID>594 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>723</ID>
<type>AA_AND2</type>
<position>298.5,-127</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>580 </input>
<output>
<ID>OUT</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>724</ID>
<type>AA_AND2</type>
<position>298.5,-131</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>725</ID>
<type>AA_AND2</type>
<position>298.5,-135</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>582 </input>
<output>
<ID>OUT</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>726</ID>
<type>AA_AND2</type>
<position>298.5,-139</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>583 </input>
<output>
<ID>OUT</ID>598 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>727</ID>
<type>AA_AND2</type>
<position>298.5,-143</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>584 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>728</ID>
<type>AA_AND2</type>
<position>298.5,-147</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>729</ID>
<type>AA_AND2</type>
<position>298.5,-151</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>586 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>730</ID>
<type>GA_LED</type>
<position>302.5,-135</position>
<input>
<ID>N_in0</ID>597 </input>
<input>
<ID>N_in1</ID>653 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>731</ID>
<type>GA_LED</type>
<position>302.5,-127</position>
<input>
<ID>N_in0</ID>596 </input>
<input>
<ID>N_in1</ID>651 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>732</ID>
<type>GA_LED</type>
<position>302.5,-131</position>
<input>
<ID>N_in0</ID>595 </input>
<input>
<ID>N_in1</ID>652 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>733</ID>
<type>GA_LED</type>
<position>302.5,-139</position>
<input>
<ID>N_in0</ID>598 </input>
<input>
<ID>N_in1</ID>654 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>734</ID>
<type>GA_LED</type>
<position>302.5,-143</position>
<input>
<ID>N_in0</ID>599 </input>
<input>
<ID>N_in1</ID>655 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>735</ID>
<type>GA_LED</type>
<position>302.5,-147</position>
<input>
<ID>N_in0</ID>600 </input>
<input>
<ID>N_in1</ID>656 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>736</ID>
<type>GA_LED</type>
<position>302.5,-151</position>
<input>
<ID>N_in0</ID>601 </input>
<input>
<ID>N_in1</ID>657 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>737</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-92</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>609 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>738</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-96</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-100</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>740</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-104</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>606 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>741</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-108</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>605 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>742</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-112</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>604 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>743</ID>
<type>AE_SMALL_INVERTER</type>
<position>293.5,-116</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>744</ID>
<type>AA_LABEL</type>
<position>265,-102</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>745</ID>
<type>AA_TOGGLE</type>
<position>276,-27</position>
<output>
<ID>OUT_0</ID>611 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>746</ID>
<type>AA_TOGGLE</type>
<position>276,-29</position>
<output>
<ID>OUT_0</ID>610 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>747</ID>
<type>AA_TOGGLE</type>
<position>276,-31</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>748</ID>
<type>AA_TOGGLE</type>
<position>276,-33</position>
<output>
<ID>OUT_0</ID>617 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>749</ID>
<type>AA_TOGGLE</type>
<position>276,-35</position>
<output>
<ID>OUT_0</ID>612 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>750</ID>
<type>AA_TOGGLE</type>
<position>276,-37</position>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>751</ID>
<type>AA_TOGGLE</type>
<position>276,-39</position>
<output>
<ID>OUT_0</ID>616 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>752</ID>
<type>AA_TOGGLE</type>
<position>276,-41</position>
<output>
<ID>OUT_0</ID>615 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>753</ID>
<type>GA_LED</type>
<position>330.5,-30</position>
<input>
<ID>N_in0</ID>626 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>754</ID>
<type>GA_LED</type>
<position>330.5,-42</position>
<input>
<ID>N_in0</ID>629 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>755</ID>
<type>GA_LED</type>
<position>330.5,-34</position>
<input>
<ID>N_in0</ID>627 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>756</ID>
<type>GA_LED</type>
<position>330.5,-38</position>
<input>
<ID>N_in0</ID>628 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>757</ID>
<type>GA_LED</type>
<position>330.5,-46</position>
<input>
<ID>N_in0</ID>630 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>758</ID>
<type>GA_LED</type>
<position>330.5,-50</position>
<input>
<ID>N_in0</ID>631 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>759</ID>
<type>GA_LED</type>
<position>330.5,-54</position>
<input>
<ID>N_in0</ID>632 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>760</ID>
<type>GA_LED</type>
<position>330.5,-58</position>
<input>
<ID>N_in0</ID>633 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>761</ID>
<type>GA_LED</type>
<position>330.5,-66.5</position>
<input>
<ID>N_in0</ID>618 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>762</ID>
<type>GA_LED</type>
<position>330.5,-78.5</position>
<input>
<ID>N_in0</ID>622 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>763</ID>
<type>GA_LED</type>
<position>330.5,-70.5</position>
<input>
<ID>N_in0</ID>619 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>764</ID>
<type>GA_LED</type>
<position>330.5,-74.5</position>
<input>
<ID>N_in0</ID>621 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>765</ID>
<type>GA_LED</type>
<position>330.5,-82.5</position>
<input>
<ID>N_in0</ID>623 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>766</ID>
<type>GA_LED</type>
<position>330.5,-86.5</position>
<input>
<ID>N_in0</ID>624 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>767</ID>
<type>GA_LED</type>
<position>330.5,-90.5</position>
<input>
<ID>N_in0</ID>625 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>768</ID>
<type>GA_LED</type>
<position>330.5,-94.5</position>
<input>
<ID>N_in0</ID>620 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>769</ID>
<type>GA_LED</type>
<position>331,-106.5</position>
<input>
<ID>N_in0</ID>650 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>770</ID>
<type>GA_LED</type>
<position>331,-118.5</position>
<input>
<ID>N_in0</ID>653 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>771</ID>
<type>GA_LED</type>
<position>331,-110.5</position>
<input>
<ID>N_in0</ID>651 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>772</ID>
<type>GA_LED</type>
<position>331,-114.5</position>
<input>
<ID>N_in0</ID>652 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>773</ID>
<type>GA_LED</type>
<position>331,-122.5</position>
<input>
<ID>N_in0</ID>654 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>774</ID>
<type>GA_LED</type>
<position>331,-126.5</position>
<input>
<ID>N_in0</ID>655 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>775</ID>
<type>GA_LED</type>
<position>331,-130.5</position>
<input>
<ID>N_in0</ID>656 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>776</ID>
<type>GA_LED</type>
<position>331,-134.5</position>
<input>
<ID>N_in0</ID>657 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>777</ID>
<type>AA_LABEL</type>
<position>338,-45</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>778</ID>
<type>AA_LABEL</type>
<position>341,-80.5</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>779</ID>
<type>AA_LABEL</type>
<position>340.5,-117.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>780</ID>
<type>AE_OR2</type>
<position>326.5,-66.5</position>
<input>
<ID>IN_0</ID>634 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>618 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>781</ID>
<type>AE_OR2</type>
<position>326.5,-70.5</position>
<input>
<ID>IN_0</ID>635 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>782</ID>
<type>AE_OR2</type>
<position>326.5,-74.5</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>644 </input>
<output>
<ID>OUT</ID>621 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>783</ID>
<type>AE_OR2</type>
<position>326.5,-78.5</position>
<input>
<ID>IN_0</ID>637 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>622 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AE_OR2</type>
<position>326.5,-82.5</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>646 </input>
<output>
<ID>OUT</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>785</ID>
<type>AE_OR2</type>
<position>326.5,-86.5</position>
<input>
<ID>IN_0</ID>639 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>624 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>AE_OR2</type>
<position>326.5,-90.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>648 </input>
<output>
<ID>OUT</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>787</ID>
<type>AE_OR2</type>
<position>326.5,-94.5</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>620 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>832</ID>
<type>AA_LABEL</type>
<position>265,-35</position>
<gparam>LABEL_TEXT ~C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1199</ID>
<type>AA_LABEL</type>
<position>60.5,-188</position>
<gparam>LABEL_TEXT Individual RGB value Selector</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1256</ID>
<type>AA_TOGGLE</type>
<position>40,-240</position>
<output>
<ID>OUT_0</ID>1021 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1257</ID>
<type>AA_LABEL</type>
<position>36.5,-239</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1258</ID>
<type>DA_FROM</type>
<position>56.5,-201</position>
<input>
<ID>IN_0</ID>1046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>1259</ID>
<type>DE_TO</type>
<position>44,-239.5</position>
<input>
<ID>IN_0</ID>1021 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>1260</ID>
<type>AA_TOGGLE</type>
<position>40,-243.5</position>
<output>
<ID>OUT_0</ID>1022 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1261</ID>
<type>DE_TO</type>
<position>44,-243.5</position>
<input>
<ID>IN_0</ID>1022 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>1262</ID>
<type>AA_TOGGLE</type>
<position>40,-245.5</position>
<output>
<ID>OUT_0</ID>1023 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1263</ID>
<type>DE_TO</type>
<position>44,-245.5</position>
<input>
<ID>IN_0</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>1264</ID>
<type>AA_TOGGLE</type>
<position>40,-247.5</position>
<output>
<ID>OUT_0</ID>1024 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1265</ID>
<type>DE_TO</type>
<position>44,-247.5</position>
<input>
<ID>IN_0</ID>1024 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>1266</ID>
<type>AA_TOGGLE</type>
<position>40,-249.5</position>
<output>
<ID>OUT_0</ID>1025 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1267</ID>
<type>DE_TO</type>
<position>44,-249.5</position>
<input>
<ID>IN_0</ID>1025 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>1268</ID>
<type>AA_TOGGLE</type>
<position>40,-251.5</position>
<output>
<ID>OUT_0</ID>1026 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1269</ID>
<type>DE_TO</type>
<position>44,-251.5</position>
<input>
<ID>IN_0</ID>1026 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>1270</ID>
<type>AA_TOGGLE</type>
<position>40,-253.5</position>
<output>
<ID>OUT_0</ID>1027 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1271</ID>
<type>DE_TO</type>
<position>44,-253.5</position>
<input>
<ID>IN_0</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>1272</ID>
<type>AA_TOGGLE</type>
<position>40,-255.5</position>
<output>
<ID>OUT_0</ID>1028 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1273</ID>
<type>DE_TO</type>
<position>44,-255.5</position>
<input>
<ID>IN_0</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>1274</ID>
<type>AA_TOGGLE</type>
<position>40,-257.5</position>
<output>
<ID>OUT_0</ID>1029 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1275</ID>
<type>DE_TO</type>
<position>44,-257.5</position>
<input>
<ID>IN_0</ID>1029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>1276</ID>
<type>DA_FROM</type>
<position>68.5,-203</position>
<input>
<ID>IN_0</ID>1030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>1277</ID>
<type>AA_LABEL</type>
<position>58,-213</position>
<gparam>LABEL_TEXT ~C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1278</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-203</position>
<input>
<ID>IN_0</ID>1030 </input>
<output>
<ID>OUT_0</ID>1038 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1279</ID>
<type>DA_FROM</type>
<position>68.5,-207</position>
<input>
<ID>IN_0</ID>1031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>1280</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-207</position>
<input>
<ID>IN_0</ID>1031 </input>
<output>
<ID>OUT_0</ID>1039 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1281</ID>
<type>DA_FROM</type>
<position>68.5,-211</position>
<input>
<ID>IN_0</ID>1032 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>1282</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-211</position>
<input>
<ID>IN_0</ID>1032 </input>
<output>
<ID>OUT_0</ID>1040 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1283</ID>
<type>DA_FROM</type>
<position>68.5,-215</position>
<input>
<ID>IN_0</ID>1033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>1284</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-215</position>
<input>
<ID>IN_0</ID>1033 </input>
<output>
<ID>OUT_0</ID>1041 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1285</ID>
<type>DA_FROM</type>
<position>68.5,-219</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>1286</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-219</position>
<input>
<ID>IN_0</ID>1034 </input>
<output>
<ID>OUT_0</ID>1042 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1287</ID>
<type>DA_FROM</type>
<position>68.5,-223</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>1288</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-223</position>
<input>
<ID>IN_0</ID>1035 </input>
<output>
<ID>OUT_0</ID>1043 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1289</ID>
<type>DA_FROM</type>
<position>68.5,-227</position>
<input>
<ID>IN_0</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>1290</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-227</position>
<input>
<ID>IN_0</ID>1036 </input>
<output>
<ID>OUT_0</ID>1044 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1291</ID>
<type>DA_FROM</type>
<position>68.5,-231</position>
<input>
<ID>IN_0</ID>1037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>1292</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-231</position>
<input>
<ID>IN_0</ID>1037 </input>
<output>
<ID>OUT_0</ID>1045 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1293</ID>
<type>AE_OR2</type>
<position>77.5,-202</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1294</ID>
<type>AE_OR2</type>
<position>77.5,-206</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1039 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1295</ID>
<type>AE_OR2</type>
<position>77.5,-210</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1040 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1296</ID>
<type>AE_OR2</type>
<position>77.5,-214</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1041 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1297</ID>
<type>AE_OR2</type>
<position>77.5,-218</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1298</ID>
<type>AE_OR2</type>
<position>77.5,-222</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1043 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1299</ID>
<type>AE_OR2</type>
<position>77.5,-226</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1044 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1300</ID>
<type>AE_OR2</type>
<position>77.5,-230</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1301</ID>
<type>AE_SMALL_INVERTER</type>
<position>60.5,-201</position>
<input>
<ID>IN_0</ID>1046 </input>
<output>
<ID>OUT_0</ID>1047 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1302</ID>
<type>DA_FROM</type>
<position>66.5,-237</position>
<input>
<ID>IN_0</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>1303</ID>
<type>DA_FROM</type>
<position>72.5,-239</position>
<input>
<ID>IN_0</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>1304</ID>
<type>AA_LABEL</type>
<position>63,-249.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1305</ID>
<type>DA_FROM</type>
<position>72.5,-243</position>
<input>
<ID>IN_0</ID>1050 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>1306</ID>
<type>DA_FROM</type>
<position>72.5,-247</position>
<input>
<ID>IN_0</ID>1051 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>1307</ID>
<type>DA_FROM</type>
<position>72.5,-251</position>
<input>
<ID>IN_0</ID>1052 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>1308</ID>
<type>DA_FROM</type>
<position>72.5,-255</position>
<input>
<ID>IN_0</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>1309</ID>
<type>DA_FROM</type>
<position>72.5,-259</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>1310</ID>
<type>DA_FROM</type>
<position>72.5,-263</position>
<input>
<ID>IN_0</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>1311</ID>
<type>DA_FROM</type>
<position>72.5,-267</position>
<input>
<ID>IN_0</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>1312</ID>
<type>AE_OR2</type>
<position>77.5,-238</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1313</ID>
<type>AE_OR2</type>
<position>77.5,-242</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1050 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1314</ID>
<type>AE_OR2</type>
<position>77.5,-246</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1051 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1315</ID>
<type>AE_OR2</type>
<position>77.5,-250</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1052 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1316</ID>
<type>AE_OR2</type>
<position>77.5,-254</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1317</ID>
<type>AE_OR2</type>
<position>77.5,-258</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1318</ID>
<type>AE_OR2</type>
<position>77.5,-262</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1319</ID>
<type>AE_OR2</type>
<position>77.5,-266</position>
<input>
<ID>IN_0</ID>1048 </input>
<input>
<ID>IN_1</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1324</ID>
<type>GA_LED</type>
<position>303.5,-508</position>
<input>
<ID>N_in0</ID>1158 </input>
<input>
<ID>N_in1</ID>167 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1325</ID>
<type>GA_LED</type>
<position>303.5,-520</position>
<input>
<ID>N_in0</ID>1161 </input>
<input>
<ID>N_in1</ID>178 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1326</ID>
<type>GA_LED</type>
<position>303.5,-512</position>
<input>
<ID>N_in0</ID>1159 </input>
<input>
<ID>N_in1</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1327</ID>
<type>GA_LED</type>
<position>303.5,-516</position>
<input>
<ID>N_in0</ID>1160 </input>
<input>
<ID>N_in1</ID>177 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1328</ID>
<type>GA_LED</type>
<position>303.5,-524</position>
<input>
<ID>N_in0</ID>1162 </input>
<input>
<ID>N_in1</ID>179 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1329</ID>
<type>GA_LED</type>
<position>303.5,-528</position>
<input>
<ID>N_in0</ID>1163 </input>
<input>
<ID>N_in1</ID>180 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1330</ID>
<type>GA_LED</type>
<position>303.5,-532</position>
<input>
<ID>N_in0</ID>1164 </input>
<input>
<ID>N_in1</ID>181 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1331</ID>
<type>GA_LED</type>
<position>303.5,-536</position>
<input>
<ID>N_in0</ID>1165 </input>
<input>
<ID>N_in1</ID>182 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1332</ID>
<type>AA_LABEL</type>
<position>310,-441</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1333</ID>
<type>AA_LABEL</type>
<position>315,-483.5</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1334</ID>
<type>AA_LABEL</type>
<position>320.5,-529.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1335</ID>
<type>AE_OR2</type>
<position>299,-468</position>
<input>
<ID>IN_0</ID>1142 </input>
<input>
<ID>IN_1</ID>1150 </input>
<output>
<ID>OUT</ID>1126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1336</ID>
<type>AE_OR2</type>
<position>299,-472</position>
<input>
<ID>IN_0</ID>1143 </input>
<input>
<ID>IN_1</ID>1151 </input>
<output>
<ID>OUT</ID>1127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1337</ID>
<type>AE_OR2</type>
<position>299,-476</position>
<input>
<ID>IN_0</ID>1144 </input>
<input>
<ID>IN_1</ID>1152 </input>
<output>
<ID>OUT</ID>1129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1338</ID>
<type>AE_OR2</type>
<position>299,-480</position>
<input>
<ID>IN_0</ID>1145 </input>
<input>
<ID>IN_1</ID>1153 </input>
<output>
<ID>OUT</ID>1130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1339</ID>
<type>AE_OR2</type>
<position>299,-484</position>
<input>
<ID>IN_0</ID>1146 </input>
<input>
<ID>IN_1</ID>1154 </input>
<output>
<ID>OUT</ID>1131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1340</ID>
<type>AE_OR2</type>
<position>299,-488</position>
<input>
<ID>IN_0</ID>1147 </input>
<input>
<ID>IN_1</ID>1155 </input>
<output>
<ID>OUT</ID>1132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1341</ID>
<type>AE_OR2</type>
<position>299,-492</position>
<input>
<ID>IN_0</ID>1148 </input>
<input>
<ID>IN_1</ID>1156 </input>
<output>
<ID>OUT</ID>1133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1342</ID>
<type>AE_OR2</type>
<position>299,-496</position>
<input>
<ID>IN_0</ID>1149 </input>
<input>
<ID>IN_1</ID>1157 </input>
<output>
<ID>OUT</ID>1128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1345</ID>
<type>GA_LED</type>
<position>275,-421</position>
<input>
<ID>N_in0</ID>1063 </input>
<input>
<ID>N_in1</ID>1134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1346</ID>
<type>AA_AND2</type>
<position>271,-421</position>
<input>
<ID>IN_0</ID>1061 </input>
<input>
<ID>IN_1</ID>1062 </input>
<output>
<ID>OUT</ID>1063 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1347</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-420</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1348</ID>
<type>AA_AND2</type>
<position>271,-425</position>
<input>
<ID>IN_0</ID>1092 </input>
<input>
<ID>IN_1</ID>1064 </input>
<output>
<ID>OUT</ID>1072 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1349</ID>
<type>AA_AND2</type>
<position>271,-429</position>
<input>
<ID>IN_0</ID>1091 </input>
<input>
<ID>IN_1</ID>1065 </input>
<output>
<ID>OUT</ID>1071 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1350</ID>
<type>AA_AND2</type>
<position>271,-433</position>
<input>
<ID>IN_0</ID>1090 </input>
<input>
<ID>IN_1</ID>1066 </input>
<output>
<ID>OUT</ID>1073 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1351</ID>
<type>AA_AND2</type>
<position>271,-437</position>
<input>
<ID>IN_0</ID>1089 </input>
<input>
<ID>IN_1</ID>1067 </input>
<output>
<ID>OUT</ID>1074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1352</ID>
<type>AA_AND2</type>
<position>271,-441</position>
<input>
<ID>IN_0</ID>1088 </input>
<input>
<ID>IN_1</ID>1068 </input>
<output>
<ID>OUT</ID>1075 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1353</ID>
<type>AA_AND2</type>
<position>271,-445</position>
<input>
<ID>IN_0</ID>1087 </input>
<input>
<ID>IN_1</ID>1069 </input>
<output>
<ID>OUT</ID>1076 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1354</ID>
<type>AA_AND2</type>
<position>271,-449</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1070 </input>
<output>
<ID>OUT</ID>1077 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1355</ID>
<type>GA_LED</type>
<position>275,-433</position>
<input>
<ID>N_in0</ID>1073 </input>
<input>
<ID>N_in1</ID>1137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1356</ID>
<type>GA_LED</type>
<position>275,-425</position>
<input>
<ID>N_in0</ID>1072 </input>
<input>
<ID>N_in1</ID>1135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1357</ID>
<type>GA_LED</type>
<position>275,-429</position>
<input>
<ID>N_in0</ID>1071 </input>
<input>
<ID>N_in1</ID>1136 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1358</ID>
<type>GA_LED</type>
<position>275,-437</position>
<input>
<ID>N_in0</ID>1074 </input>
<input>
<ID>N_in1</ID>1138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1359</ID>
<type>GA_LED</type>
<position>275,-441</position>
<input>
<ID>N_in0</ID>1075 </input>
<input>
<ID>N_in1</ID>1139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1360</ID>
<type>GA_LED</type>
<position>275,-445</position>
<input>
<ID>N_in0</ID>1076 </input>
<input>
<ID>N_in1</ID>1140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1361</ID>
<type>GA_LED</type>
<position>275,-449</position>
<input>
<ID>N_in0</ID>1077 </input>
<input>
<ID>N_in1</ID>1141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1362</ID>
<type>GA_LED</type>
<position>275,-455</position>
<input>
<ID>N_in0</ID>1078 </input>
<input>
<ID>N_in1</ID>1142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1363</ID>
<type>AA_AND2</type>
<position>271,-455</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1062 </input>
<output>
<ID>OUT</ID>1078 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1364</ID>
<type>AA_AND2</type>
<position>271,-459</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1064 </input>
<output>
<ID>OUT</ID>1080 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1365</ID>
<type>AA_AND2</type>
<position>271,-463</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1065 </input>
<output>
<ID>OUT</ID>1079 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1366</ID>
<type>AA_AND2</type>
<position>271,-467</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1066 </input>
<output>
<ID>OUT</ID>1081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1367</ID>
<type>AA_AND2</type>
<position>271,-471</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1067 </input>
<output>
<ID>OUT</ID>1082 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1368</ID>
<type>AA_AND2</type>
<position>271,-475</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1068 </input>
<output>
<ID>OUT</ID>1083 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1369</ID>
<type>AA_AND2</type>
<position>271,-479</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1069 </input>
<output>
<ID>OUT</ID>1084 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1370</ID>
<type>AA_AND2</type>
<position>271,-483</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1070 </input>
<output>
<ID>OUT</ID>1085 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1371</ID>
<type>GA_LED</type>
<position>275,-467</position>
<input>
<ID>N_in0</ID>1081 </input>
<input>
<ID>N_in1</ID>1145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1372</ID>
<type>GA_LED</type>
<position>275,-459</position>
<input>
<ID>N_in0</ID>1080 </input>
<input>
<ID>N_in1</ID>1143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1373</ID>
<type>GA_LED</type>
<position>275,-463</position>
<input>
<ID>N_in0</ID>1079 </input>
<input>
<ID>N_in1</ID>1144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1374</ID>
<type>GA_LED</type>
<position>275,-471</position>
<input>
<ID>N_in0</ID>1082 </input>
<input>
<ID>N_in1</ID>1146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1375</ID>
<type>GA_LED</type>
<position>275,-475</position>
<input>
<ID>N_in0</ID>1083 </input>
<input>
<ID>N_in1</ID>1147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1376</ID>
<type>GA_LED</type>
<position>275,-479</position>
<input>
<ID>N_in0</ID>1084 </input>
<input>
<ID>N_in1</ID>1148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1377</ID>
<type>GA_LED</type>
<position>275,-483</position>
<input>
<ID>N_in0</ID>1085 </input>
<input>
<ID>N_in1</ID>1149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1378</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-424</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1092 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1379</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-428</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1091 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1380</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-432</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1090 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1381</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-436</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1089 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1382</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-440</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1088 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1383</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-444</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1087 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1384</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-448</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1086 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1386</ID>
<type>GA_LED</type>
<position>275,-490.5</position>
<input>
<ID>N_in0</ID>1095 </input>
<input>
<ID>N_in1</ID>1150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1387</ID>
<type>AA_AND2</type>
<position>271,-490.5</position>
<input>
<ID>IN_0</ID>1093 </input>
<input>
<ID>IN_1</ID>1094 </input>
<output>
<ID>OUT</ID>1095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1388</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-489.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1093 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1389</ID>
<type>AA_AND2</type>
<position>271,-494.5</position>
<input>
<ID>IN_0</ID>1125 </input>
<input>
<ID>IN_1</ID>1096 </input>
<output>
<ID>OUT</ID>1104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1390</ID>
<type>AA_AND2</type>
<position>271,-498.5</position>
<input>
<ID>IN_0</ID>1124 </input>
<input>
<ID>IN_1</ID>1097 </input>
<output>
<ID>OUT</ID>1103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1391</ID>
<type>AA_AND2</type>
<position>271,-502.5</position>
<input>
<ID>IN_0</ID>1123 </input>
<input>
<ID>IN_1</ID>1098 </input>
<output>
<ID>OUT</ID>1105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1392</ID>
<type>AA_AND2</type>
<position>271,-506.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<input>
<ID>IN_1</ID>1099 </input>
<output>
<ID>OUT</ID>1106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1393</ID>
<type>AA_AND2</type>
<position>271,-510.5</position>
<input>
<ID>IN_0</ID>1121 </input>
<input>
<ID>IN_1</ID>1100 </input>
<output>
<ID>OUT</ID>1107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1394</ID>
<type>AA_AND2</type>
<position>271,-514.5</position>
<input>
<ID>IN_0</ID>1120 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1395</ID>
<type>AA_AND2</type>
<position>271,-518.5</position>
<input>
<ID>IN_0</ID>1118 </input>
<input>
<ID>IN_1</ID>1102 </input>
<output>
<ID>OUT</ID>1109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1396</ID>
<type>GA_LED</type>
<position>275,-502.5</position>
<input>
<ID>N_in0</ID>1105 </input>
<input>
<ID>N_in1</ID>1153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1397</ID>
<type>GA_LED</type>
<position>275,-494.5</position>
<input>
<ID>N_in0</ID>1104 </input>
<input>
<ID>N_in1</ID>1151 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1398</ID>
<type>GA_LED</type>
<position>275,-498.5</position>
<input>
<ID>N_in0</ID>1103 </input>
<input>
<ID>N_in1</ID>1152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1399</ID>
<type>GA_LED</type>
<position>275,-506.5</position>
<input>
<ID>N_in0</ID>1106 </input>
<input>
<ID>N_in1</ID>1154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1400</ID>
<type>GA_LED</type>
<position>275,-510.5</position>
<input>
<ID>N_in0</ID>1107 </input>
<input>
<ID>N_in1</ID>1155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1401</ID>
<type>GA_LED</type>
<position>275,-514.5</position>
<input>
<ID>N_in0</ID>1108 </input>
<input>
<ID>N_in1</ID>1156 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1402</ID>
<type>GA_LED</type>
<position>275,-518.5</position>
<input>
<ID>N_in0</ID>1109 </input>
<input>
<ID>N_in1</ID>1157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1403</ID>
<type>GA_LED</type>
<position>275,-524.5</position>
<input>
<ID>N_in0</ID>1110 </input>
<input>
<ID>N_in1</ID>1158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1404</ID>
<type>AA_AND2</type>
<position>271,-524.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1094 </input>
<output>
<ID>OUT</ID>1110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1405</ID>
<type>AA_AND2</type>
<position>271,-528.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1096 </input>
<output>
<ID>OUT</ID>1112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1406</ID>
<type>AA_AND2</type>
<position>271,-532.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1097 </input>
<output>
<ID>OUT</ID>1111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1407</ID>
<type>AA_AND2</type>
<position>271,-536.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1098 </input>
<output>
<ID>OUT</ID>1113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1408</ID>
<type>AA_AND2</type>
<position>271,-540.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1099 </input>
<output>
<ID>OUT</ID>1114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1409</ID>
<type>AA_AND2</type>
<position>271,-544.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1100 </input>
<output>
<ID>OUT</ID>1115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1410</ID>
<type>AA_AND2</type>
<position>271,-548.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1411</ID>
<type>AA_AND2</type>
<position>271,-552.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1102 </input>
<output>
<ID>OUT</ID>1117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1412</ID>
<type>GA_LED</type>
<position>275,-536.5</position>
<input>
<ID>N_in0</ID>1113 </input>
<input>
<ID>N_in1</ID>1161 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1413</ID>
<type>GA_LED</type>
<position>275,-528.5</position>
<input>
<ID>N_in0</ID>1112 </input>
<input>
<ID>N_in1</ID>1159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1414</ID>
<type>GA_LED</type>
<position>275,-532.5</position>
<input>
<ID>N_in0</ID>1111 </input>
<input>
<ID>N_in1</ID>1160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1415</ID>
<type>GA_LED</type>
<position>275,-540.5</position>
<input>
<ID>N_in0</ID>1114 </input>
<input>
<ID>N_in1</ID>1162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1416</ID>
<type>GA_LED</type>
<position>275,-544.5</position>
<input>
<ID>N_in0</ID>1115 </input>
<input>
<ID>N_in1</ID>1163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1417</ID>
<type>GA_LED</type>
<position>275,-548.5</position>
<input>
<ID>N_in0</ID>1116 </input>
<input>
<ID>N_in1</ID>1164 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1418</ID>
<type>GA_LED</type>
<position>275,-552.5</position>
<input>
<ID>N_in0</ID>1117 </input>
<input>
<ID>N_in1</ID>1165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1419</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-493.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1125 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1420</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-497.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1124 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1421</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-501.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1123 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1422</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-505.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1122 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1423</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-509.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1121 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1424</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-513.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1120 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1425</ID>
<type>AE_SMALL_INVERTER</type>
<position>266,-517.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<output>
<ID>OUT_0</ID>1118 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1426</ID>
<type>GA_LED</type>
<position>303,-431.5</position>
<input>
<ID>N_in0</ID>1134 </input>
<input>
<ID>N_in1</ID>151 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1427</ID>
<type>GA_LED</type>
<position>303,-443.5</position>
<input>
<ID>N_in0</ID>1137 </input>
<input>
<ID>N_in1</ID>154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1428</ID>
<type>GA_LED</type>
<position>303,-435.5</position>
<input>
<ID>N_in0</ID>1135 </input>
<input>
<ID>N_in1</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1429</ID>
<type>GA_LED</type>
<position>303,-439.5</position>
<input>
<ID>N_in0</ID>1136 </input>
<input>
<ID>N_in1</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1430</ID>
<type>GA_LED</type>
<position>303,-447.5</position>
<input>
<ID>N_in0</ID>1138 </input>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1431</ID>
<type>GA_LED</type>
<position>303,-451.5</position>
<input>
<ID>N_in0</ID>1139 </input>
<input>
<ID>N_in1</ID>156 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1432</ID>
<type>GA_LED</type>
<position>303,-455.5</position>
<input>
<ID>N_in0</ID>1140 </input>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1433</ID>
<type>GA_LED</type>
<position>303,-459.5</position>
<input>
<ID>N_in0</ID>1141 </input>
<input>
<ID>N_in1</ID>158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1434</ID>
<type>GA_LED</type>
<position>303,-468</position>
<input>
<ID>N_in0</ID>1126 </input>
<input>
<ID>N_in1</ID>159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1435</ID>
<type>GA_LED</type>
<position>303,-480</position>
<input>
<ID>N_in0</ID>1130 </input>
<input>
<ID>N_in1</ID>162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1436</ID>
<type>GA_LED</type>
<position>303,-472</position>
<input>
<ID>N_in0</ID>1127 </input>
<input>
<ID>N_in1</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1437</ID>
<type>GA_LED</type>
<position>303,-476</position>
<input>
<ID>N_in0</ID>1129 </input>
<input>
<ID>N_in1</ID>161 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1438</ID>
<type>GA_LED</type>
<position>303,-484</position>
<input>
<ID>N_in0</ID>1131 </input>
<input>
<ID>N_in1</ID>163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1439</ID>
<type>GA_LED</type>
<position>303,-488</position>
<input>
<ID>N_in0</ID>1132 </input>
<input>
<ID>N_in1</ID>164 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1440</ID>
<type>GA_LED</type>
<position>303,-492</position>
<input>
<ID>N_in0</ID>1133 </input>
<input>
<ID>N_in1</ID>165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1441</ID>
<type>GA_LED</type>
<position>303,-496</position>
<input>
<ID>N_in0</ID>1128 </input>
<input>
<ID>N_in1</ID>166 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1463</ID>
<type>AA_LABEL</type>
<position>226.5,-433</position>
<gparam>LABEL_TEXT ~C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1464</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-423</position>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>1183 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1466</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-427</position>
<input>
<ID>IN_0</ID>149 </input>
<output>
<ID>OUT_0</ID>1184 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1468</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-431</position>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>1185 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1470</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-435</position>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT_0</ID>1186 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1472</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-439</position>
<input>
<ID>IN_0</ID>146 </input>
<output>
<ID>OUT_0</ID>1187 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1474</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-443</position>
<input>
<ID>IN_0</ID>145 </input>
<output>
<ID>OUT_0</ID>1188 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1476</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-447</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>1189 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1478</ID>
<type>AE_SMALL_INVERTER</type>
<position>241,-451</position>
<input>
<ID>IN_0</ID>143 </input>
<output>
<ID>OUT_0</ID>1190 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1479</ID>
<type>AE_OR2</type>
<position>246,-422</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1183 </input>
<output>
<ID>OUT</ID>1062 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1480</ID>
<type>AE_OR2</type>
<position>246,-426</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1184 </input>
<output>
<ID>OUT</ID>1064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1481</ID>
<type>AE_OR2</type>
<position>246,-430</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1185 </input>
<output>
<ID>OUT</ID>1065 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1482</ID>
<type>AE_OR2</type>
<position>246,-434</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1186 </input>
<output>
<ID>OUT</ID>1066 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1483</ID>
<type>AE_OR2</type>
<position>246,-438</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1187 </input>
<output>
<ID>OUT</ID>1067 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1484</ID>
<type>AE_OR2</type>
<position>246,-442</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1188 </input>
<output>
<ID>OUT</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1485</ID>
<type>AE_OR2</type>
<position>246,-446</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1189 </input>
<output>
<ID>OUT</ID>1069 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1486</ID>
<type>AE_OR2</type>
<position>246,-450</position>
<input>
<ID>IN_0</ID>1192 </input>
<input>
<ID>IN_1</ID>1190 </input>
<output>
<ID>OUT</ID>1070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1487</ID>
<type>AE_SMALL_INVERTER</type>
<position>229,-421</position>
<input>
<ID>IN_0</ID>1193 </input>
<output>
<ID>OUT_0</ID>1192 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1490</ID>
<type>AA_LABEL</type>
<position>231,-503</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1498</ID>
<type>AE_OR2</type>
<position>245.5,-491.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>1094 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1499</ID>
<type>AE_OR2</type>
<position>245.5,-495.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>1096 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1500</ID>
<type>AE_OR2</type>
<position>245.5,-499.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>1097 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1501</ID>
<type>AE_OR2</type>
<position>245.5,-503.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>1098 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1502</ID>
<type>AE_OR2</type>
<position>245.5,-507.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>1099 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1503</ID>
<type>AE_OR2</type>
<position>245.5,-511.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>1100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1504</ID>
<type>AE_OR2</type>
<position>245.5,-515.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>1101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1505</ID>
<type>AE_OR2</type>
<position>245.5,-519.5</position>
<input>
<ID>IN_0</ID>1193 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>1102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1506</ID>
<type>AE_REGISTER8</type>
<position>322,-447.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>154 </input>
<input>
<ID>IN_4</ID>155 </input>
<input>
<ID>IN_5</ID>156 </input>
<input>
<ID>IN_6</ID>157 </input>
<input>
<ID>IN_7</ID>158 </input>
<input>
<ID>clock</ID>1203 </input>
<input>
<ID>load</ID>1204 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1507</ID>
<type>AE_REGISTER8</type>
<position>326,-521</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<input>
<ID>IN_2</ID>177 </input>
<input>
<ID>IN_3</ID>178 </input>
<input>
<ID>IN_4</ID>179 </input>
<input>
<ID>IN_5</ID>180 </input>
<input>
<ID>IN_6</ID>181 </input>
<input>
<ID>IN_7</ID>182 </input>
<input>
<ID>clock</ID>1202 </input>
<input>
<ID>load</ID>1207 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1508</ID>
<type>BB_CLOCK</type>
<position>318.5,-533</position>
<output>
<ID>CLK</ID>1202 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1509</ID>
<type>BB_CLOCK</type>
<position>316,-455.5</position>
<output>
<ID>CLK</ID>1203 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1510</ID>
<type>AA_TOGGLE</type>
<position>318.5,-440.5</position>
<output>
<ID>OUT_0</ID>1204 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1511</ID>
<type>AE_REGISTER8</type>
<position>324,-479.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>160 </input>
<input>
<ID>IN_2</ID>161 </input>
<input>
<ID>IN_3</ID>162 </input>
<input>
<ID>IN_4</ID>163 </input>
<input>
<ID>IN_5</ID>164 </input>
<input>
<ID>IN_6</ID>165 </input>
<input>
<ID>IN_7</ID>166 </input>
<input>
<ID>clock</ID>1205 </input>
<input>
<ID>load</ID>1206 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1512</ID>
<type>BB_CLOCK</type>
<position>317,-489.5</position>
<output>
<ID>CLK</ID>1205 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1513</ID>
<type>AA_TOGGLE</type>
<position>320.5,-472</position>
<output>
<ID>OUT_0</ID>1206 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1514</ID>
<type>AA_TOGGLE</type>
<position>321.5,-511</position>
<output>
<ID>OUT_0</ID>1207 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1515</ID>
<type>BE_JKFF_LOW</type>
<position>113,72</position>
<input>
<ID>J</ID>1208 </input>
<input>
<ID>K</ID>1208 </input>
<input>
<ID>clock</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1517</ID>
<type>AA_LABEL</type>
<position>90.5,78.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1519</ID>
<type>AA_TOGGLE</type>
<position>94.5,69</position>
<output>
<ID>OUT_0</ID>322 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1521</ID>
<type>AE_REGISTER8</type>
<position>99.5,59</position>
<output>
<ID>carry_out</ID>1208 </output>
<input>
<ID>clock</ID>312 </input>
<input>
<ID>count_enable</ID>1210 </input>
<input>
<ID>count_up</ID>1212 </input>
<input>
<ID>load</ID>322 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1531</ID>
<type>BE_JKFF_LOW</type>
<position>99,78</position>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1532</ID>
<type>BE_JKFF_LOW</type>
<position>99,87.5</position>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>157.5,-502,199.5,-502</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>162 5</intersection>
<intersection>173.5 8</intersection>
<intersection>199.5 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>162,-502,162,-489</points>
<connection>
<GID>253</GID>
<name>clear</name></connection>
<intersection>-502 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>199.5,-502,199.5,-472.5</points>
<connection>
<GID>232</GID>
<name>clear</name></connection>
<intersection>-502 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>173.5,-502,173.5,-472.5</points>
<intersection>-502 2</intersection>
<intersection>-472.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>173.5,-472.5,176.5,-472.5</points>
<connection>
<GID>231</GID>
<name>clear</name></connection>
<intersection>173.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,125.5,78,137.5</points>
<intersection>125.5 4</intersection>
<intersection>129.5 1</intersection>
<intersection>137.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,129.5,79,129.5</points>
<connection>
<GID>5</GID>
<name>J</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>78,125.5,79,125.5</points>
<connection>
<GID>5</GID>
<name>K</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>77,137.5,78,137.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,117.5,98,117.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>79 4</intersection>
<intersection>98 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>98,117.5,98,127.5</points>
<intersection>117.5 1</intersection>
<intersection>127.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>79,117.5,79,127.5</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>117.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>98,127.5,102,127.5</points>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<intersection>98 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,120,85,120</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-19,43.5,-19</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-25.5,32.5,-12</points>
<intersection>-25.5 4</intersection>
<intersection>-19 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-19,36,-19</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-12,32.5,-12</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-25.5,43,-25.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-27.5,43,-27.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-27.5,40,-21</points>
<intersection>-27.5 1</intersection>
<intersection>-21 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>40,-21,43.5,-21</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>40 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-20,56,-20</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-26.5,56,-26.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,120,74.5,134.5</points>
<intersection>120 1</intersection>
<intersection>127.5 2</intersection>
<intersection>134.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,120,80.5,120</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,127.5,74.5,127.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,134.5,86,134.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,122,85,125.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>nQ</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,129.5,85,139.5</points>
<connection>
<GID>5</GID>
<name>Q</name></connection>
<connection>
<GID>56</GID>
<name>N_in2</name></connection>
<intersection>132.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>85,132.5,86,132.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,130.5,92,133.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,121,92,128.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>121 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>91,121,92,121</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-23,118.5,-23</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,125.5,99.5,129.5</points>
<intersection>125.5 3</intersection>
<intersection>129.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,129.5,102,129.5</points>
<connection>
<GID>9</GID>
<name>J</name></connection>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99.5,125.5,102,125.5</points>
<connection>
<GID>9</GID>
<name>K</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-31.5,108,-31.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,-59,108,-25</points>
<intersection>-59 19</intersection>
<intersection>-31.5 1</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>108,-25,118.5,-25</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>108 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>108,-59,118.5,-59</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>108 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>124.5,-24,124.5,-24</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,129.5,108,138.5</points>
<connection>
<GID>9</GID>
<name>Q</name></connection>
<connection>
<GID>58</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-63,108.5,-29</points>
<intersection>-63 3</intersection>
<intersection>-33.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-29,118.5,-29</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-33.5,108.5,-33.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108.5,-63,118.5,-63</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-67,109,-33</points>
<intersection>-67 3</intersection>
<intersection>-35.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-33,118.5,-33</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-35.5,109,-35.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>109,-67,118.5,-67</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>109 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-37.5,109.5,-37.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>109.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>109.5,-71,109.5,-37</points>
<intersection>-71 5</intersection>
<intersection>-37.5 1</intersection>
<intersection>-37 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>109.5,-71,118.5,-71</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>109.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>109.5,-37,118.5,-37</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>109.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-39.5,110,-39.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-75,110,-39.5</points>
<intersection>-75 4</intersection>
<intersection>-41 8</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>110,-75,118.5,-75</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>110 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>110,-41,118.5,-41</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>110 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-41.5,110.5,-41.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>110.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110.5,-79,110.5,-41.5</points>
<intersection>-79 4</intersection>
<intersection>-45 8</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>110.5,-79,118.5,-79</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>110.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>110.5,-45,118.5,-45</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>110.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-49,109,-43.5</points>
<intersection>-49 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109,-49,118.5,-49</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>109 0</intersection>
<intersection>111 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-43.5,109,-43.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>109 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-83,111,-49</points>
<intersection>-83 4</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>111,-83,118.5,-83</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>111 3</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-45.5,111.5,-45.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>111.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111.5,-87,111.5,-45.5</points>
<intersection>-87 4</intersection>
<intersection>-53 5</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>111.5,-87,118.5,-87</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>111.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>111.5,-53,118.5,-53</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>111.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230,93,230,105</points>
<intersection>93 4</intersection>
<intersection>97 1</intersection>
<intersection>105 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230,97,231,97</points>
<connection>
<GID>100</GID>
<name>J</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>230,93,231,93</points>
<connection>
<GID>100</GID>
<name>K</name></connection>
<intersection>230 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>229,105,230,105</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>230 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,85.5,253,85.5</points>
<connection>
<GID>226</GID>
<name>carry_out</name></connection>
<intersection>228 6</intersection>
<intersection>253 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>228,85.5,228,95</points>
<intersection>85.5 1</intersection>
<intersection>95 8</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>253,85.5,253,95</points>
<intersection>85.5 1</intersection>
<intersection>95 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>228,95,231,95</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<intersection>228 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>253,95,254,95</points>
<connection>
<GID>101</GID>
<name>clock</name></connection>
<intersection>253 7</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,87.5,237,87.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-203.5,195,-203.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,89.5,237,93</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>nQ</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-32,124.5,-32</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-28,124.5,-28</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<connection>
<GID>61</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-36,124.5,-36</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>60</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-40,124.5,-40</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-44,124.5,-44</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>64</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-48,124.5,-48</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-52,124.5,-52</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237,97,237,107</points>
<connection>
<GID>100</GID>
<name>Q</name></connection>
<connection>
<GID>201</GID>
<name>N_in2</name></connection>
<intersection>100 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>237,100,238,100</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>237 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>124.5,-58,124.5,-58</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-66,124.5,-66</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<connection>
<GID>78</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-62,124.5,-62</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-70,124.5,-70</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-74,124.5,-74</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-78,124.5,-78</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-82,124.5,-82</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<connection>
<GID>81</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-86,124.5,-86</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-51,118.5,-51</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-85,107.5,-16</points>
<intersection>-85 18</intersection>
<intersection>-81 17</intersection>
<intersection>-77 16</intersection>
<intersection>-73 15</intersection>
<intersection>-69 14</intersection>
<intersection>-65 13</intersection>
<intersection>-61 12</intersection>
<intersection>-57 11</intersection>
<intersection>-51 2</intersection>
<intersection>-47 9</intersection>
<intersection>-43 8</intersection>
<intersection>-39 7</intersection>
<intersection>-35 6</intersection>
<intersection>-31 5</intersection>
<intersection>-27 4</intersection>
<intersection>-23 3</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-16,107.5,-16</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107.5,-51,114.5,-51</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-23,114.5,-23</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>107.5,-27,114.5,-27</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>107.5,-31,114.5,-31</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>107.5,-35,114.5,-35</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>107.5,-39,114.5,-39</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>107.5,-43,114.5,-43</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>107.5,-47,114.5,-47</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>107.5,-57,118.5,-57</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>107.5,-61,118.5,-61</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>107.5,-65,118.5,-65</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>107.5,-69,118.5,-69</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>107.5,-73,118.5,-73</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>107.5,-77,118.5,-77</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>107.5,-81,118.5,-81</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>107.5,-85,118.5,-85</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-47,118.5,-47</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-43,118.5,-43</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-39,118.5,-39</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-35,118.5,-35</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-31,118.5,-31</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>118.5,-27,118.5,-27</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-21,208.5,-21</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>198,-57,198,-23</points>
<intersection>-57 19</intersection>
<intersection>-29.5 23</intersection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>198,-23,208.5,-23</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>198 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>198,-57,208.5,-57</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>198 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>195,-29.5,198,-29.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>198 3</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>214.5,-22,214.5,-22</points>
<connection>
<GID>95</GID>
<name>N_in0</name></connection>
<connection>
<GID>96</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-61,198.5,-27</points>
<intersection>-61 3</intersection>
<intersection>-31.5 6</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198.5,-27,208.5,-27</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-61,208.5,-61</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>195,-31.5,198.5,-31.5</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-65,199,-31</points>
<intersection>-65 3</intersection>
<intersection>-33.5 6</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-31,208.5,-31</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>199,-65,208.5,-65</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>195,-33.5,199,-33.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>199 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>199.5,-69,199.5,-35</points>
<intersection>-69 5</intersection>
<intersection>-35.5 11</intersection>
<intersection>-35 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>199.5,-69,208.5,-69</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>199.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>199.5,-35,208.5,-35</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>199.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>195,-35.5,199.5,-35.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>199.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>200,-73,200,-37.5</points>
<intersection>-73 4</intersection>
<intersection>-39 8</intersection>
<intersection>-37.5 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>200,-73,208.5,-73</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>200 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200,-39,208.5,-39</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>200 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>195,-37.5,200,-37.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>200 3</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-39.5,208.5,-39.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>200.5 3</intersection>
<intersection>208.5 11</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>200.5,-77,200.5,-39.5</points>
<intersection>-77 4</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>200.5,-77,208.5,-77</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>200.5 3</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>208.5,-43,208.5,-39.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>201,-47,208.5,-47</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>201 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201,-81,201,-41.5</points>
<intersection>-81 4</intersection>
<intersection>-47 1</intersection>
<intersection>-41.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>201,-81,208.5,-81</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>201 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>195,-41.5,201,-41.5</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>201 3</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>201.5,-85,201.5,-43.5</points>
<intersection>-85 4</intersection>
<intersection>-51 5</intersection>
<intersection>-43.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>201.5,-85,208.5,-85</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>201.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>201.5,-51,208.5,-51</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>201.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>195,-43.5,201.5,-43.5</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>201.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-30,214.5,-30</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-26,214.5,-26</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>113</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-34,214.5,-34</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-38,214.5,-38</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-42,214.5,-42</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-46,214.5,-46</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<connection>
<GID>117</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-50,214.5,-50</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>214.5,-56,214.5,-56</points>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-64,214.5,-64</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<connection>
<GID>130</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-60,214.5,-60</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-68,214.5,-68</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-72,214.5,-72</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-76,214.5,-76</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>132</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-80,214.5,-80</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<connection>
<GID>133</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-84,214.5,-84</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-49,208.5,-49</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,98,244,101</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-45,208.5,-45</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-41,208.5,-41</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-37,208.5,-37</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-33,208.5,-33</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-29,208.5,-29</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-25,208.5,-25</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-90.5,208.5,-90.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-99,198,-99</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>198 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>198,-126.5,198,-92.5</points>
<intersection>-126.5 19</intersection>
<intersection>-99 1</intersection>
<intersection>-92.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>198,-92.5,208.5,-92.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>198 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>198,-126.5,208.5,-126.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>198 3</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>214.5,-91.5,214.5,-91.5</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<connection>
<GID>146</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198.5,-130.5,198.5,-96.5</points>
<intersection>-130.5 3</intersection>
<intersection>-101 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198.5,-96.5,208.5,-96.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-101,198.5,-101</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>198.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>198.5,-130.5,208.5,-130.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-134.5,199,-100.5</points>
<intersection>-134.5 3</intersection>
<intersection>-103 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-100.5,208.5,-100.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-103,199,-103</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>199,-134.5,208.5,-134.5</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-105,199.5,-105</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>199.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>199.5,-138.5,199.5,-104.5</points>
<intersection>-138.5 5</intersection>
<intersection>-105 1</intersection>
<intersection>-104.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>199.5,-138.5,208.5,-138.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>199.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>199.5,-104.5,208.5,-104.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>199.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-107,200,-107</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>200 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>200,-142.5,200,-107</points>
<intersection>-142.5 4</intersection>
<intersection>-108.5 8</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>200,-142.5,208.5,-142.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>200 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200,-108.5,208.5,-108.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>200 3</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-109,200.5,-109</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>200.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>200.5,-146.5,200.5,-109</points>
<intersection>-146.5 4</intersection>
<intersection>-112.5 8</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>200.5,-146.5,208.5,-146.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>200.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,-112.5,208.5,-112.5</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>200.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-116.5,199,-111</points>
<intersection>-116.5 1</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-116.5,208.5,-116.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection>
<intersection>201 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-111,199,-111</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>199 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201,-150.5,201,-116.5</points>
<intersection>-150.5 4</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>201,-150.5,208.5,-150.5</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>201 3</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194.5,-113,201.5,-113</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>201.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201.5,-154.5,201.5,-113</points>
<intersection>-154.5 4</intersection>
<intersection>-120.5 5</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>201.5,-154.5,208.5,-154.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>201.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>201.5,-120.5,208.5,-120.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>201.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-99.5,214.5,-99.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<connection>
<GID>164</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-95.5,214.5,-95.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<connection>
<GID>163</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-103.5,214.5,-103.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-107.5,214.5,-107.5</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-111.5,214.5,-111.5</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<connection>
<GID>166</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-115.5,214.5,-115.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<connection>
<GID>167</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-119.5,214.5,-119.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<connection>
<GID>168</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>214.5,-125.5,214.5,-125.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<connection>
<GID>170</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-133.5,214.5,-133.5</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<connection>
<GID>180</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-129.5,214.5,-129.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<connection>
<GID>179</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-137.5,214.5,-137.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-141.5,214.5,-141.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<connection>
<GID>181</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-145.5,214.5,-145.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>182</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-149.5,214.5,-149.5</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>183</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-153.5,214.5,-153.5</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<connection>
<GID>184</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-118.5,208.5,-118.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-152.5,197.5,-14</points>
<intersection>-152.5 18</intersection>
<intersection>-148.5 17</intersection>
<intersection>-144.5 16</intersection>
<intersection>-140.5 15</intersection>
<intersection>-136.5 14</intersection>
<intersection>-132.5 13</intersection>
<intersection>-128.5 12</intersection>
<intersection>-124.5 11</intersection>
<intersection>-118.5 2</intersection>
<intersection>-114.5 9</intersection>
<intersection>-110.5 8</intersection>
<intersection>-106.5 7</intersection>
<intersection>-102.5 6</intersection>
<intersection>-98.5 5</intersection>
<intersection>-94.5 4</intersection>
<intersection>-90.5 3</intersection>
<intersection>-83 38</intersection>
<intersection>-79 37</intersection>
<intersection>-75 36</intersection>
<intersection>-71 35</intersection>
<intersection>-67 34</intersection>
<intersection>-63 33</intersection>
<intersection>-59 32</intersection>
<intersection>-55 31</intersection>
<intersection>-49 22</intersection>
<intersection>-45 29</intersection>
<intersection>-41 28</intersection>
<intersection>-37 27</intersection>
<intersection>-33 26</intersection>
<intersection>-29 25</intersection>
<intersection>-25 24</intersection>
<intersection>-21 23</intersection>
<intersection>-14 21</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>197.5,-118.5,204.5,-118.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>197.5,-90.5,204.5,-90.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>197.5,-94.5,204.5,-94.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>197.5,-98.5,204.5,-98.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>197.5,-102.5,204.5,-102.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>197.5,-106.5,204.5,-106.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>197.5,-110.5,204.5,-110.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>197.5,-114.5,204.5,-114.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>197.5,-124.5,208.5,-124.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>197.5,-128.5,208.5,-128.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>197.5,-132.5,208.5,-132.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>197.5,-136.5,208.5,-136.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>197.5,-140.5,208.5,-140.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>197.5,-144.5,208.5,-144.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>197.5,-148.5,208.5,-148.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>197.5,-152.5,208.5,-152.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>185,-14,197.5,-14</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>197.5,-49,204.5,-49</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>197.5,-21,204.5,-21</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>197.5,-25,204.5,-25</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>197.5,-29,204.5,-29</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>197.5,-33,204.5,-33</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>197.5,-37,204.5,-37</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>197.5,-41,204.5,-41</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>197.5,-45,204.5,-45</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>197.5,-55,208.5,-55</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>197.5,-59,208.5,-59</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>197.5,-63,208.5,-63</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>197.5,-67,208.5,-67</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>197.5,-71,208.5,-71</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>197.5,-75,208.5,-75</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>197.5,-79,208.5,-79</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>197.5,-83,208.5,-83</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-114.5,208.5,-114.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-110.5,208.5,-110.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-106.5,208.5,-106.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-102.5,208.5,-102.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-98.5,208.5,-98.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208.5,-94.5,208.5,-94.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,88.5,244,96</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>88.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>243,88.5,244,88.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,93,251.5,97</points>
<intersection>93 3</intersection>
<intersection>97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,97,254,97</points>
<connection>
<GID>101</GID>
<name>J</name></connection>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>251.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>251.5,93,254,93</points>
<connection>
<GID>101</GID>
<name>K</name></connection>
<intersection>251.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>260,97,260,106</points>
<connection>
<GID>101</GID>
<name>Q</name></connection>
<connection>
<GID>202</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,69.5,217.5,74.5</points>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<intersection>69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,69.5,217.5,69.5</points>
<intersection>192.5 2</intersection>
<intersection>217.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>192.5,69.5,192.5,79</points>
<intersection>69.5 1</intersection>
<intersection>79 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>188,79,192.5,79</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>192.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>217,87,217,89.5</points>
<intersection>87 34</intersection>
<intersection>89.5 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>215.5,89.5,218.5,89.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>217 5</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>217,87,217.5,87</points>
<intersection>217 5</intersection>
<intersection>217.5 35</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>217.5,85.5,217.5,87</points>
<connection>
<GID>226</GID>
<name>load</name></connection>
<intersection>87 34</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>184.5,-239.5,184.5,-205.5</points>
<intersection>-239.5 19</intersection>
<intersection>-205.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>176,-205.5,195,-205.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>184.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>184.5,-239.5,195,-239.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>184.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,85.5,218.5,85.5</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<connection>
<GID>226</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,85.5,219.5,92</points>
<connection>
<GID>226</GID>
<name>count_up</name></connection>
<intersection>92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,92,219.5,92</points>
<intersection>195.5 2</intersection>
<intersection>219.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>195.5,75,195.5,95</points>
<intersection>75 3</intersection>
<intersection>92 1</intersection>
<intersection>95 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>188,75,195.5,75</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>195.5 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>225.5,87.5,225.5,102</points>
<intersection>87.5 6</intersection>
<intersection>95 7</intersection>
<intersection>102 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>225.5,87.5,232.5,87.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>225.5 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>195.5,95,225.5,95</points>
<intersection>195.5 2</intersection>
<intersection>225.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>225.5,102,238,102</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>225.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-470.5,172.5,-458.5</points>
<intersection>-470.5 4</intersection>
<intersection>-466.5 1</intersection>
<intersection>-458.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,-466.5,173.5,-466.5</points>
<connection>
<GID>231</GID>
<name>J</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>172.5,-470.5,173.5,-470.5</points>
<connection>
<GID>231</GID>
<name>K</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>171.5,-458.5,172.5,-458.5</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163,-478,195.5,-478</points>
<connection>
<GID>253</GID>
<name>carry_out</name></connection>
<intersection>170.5 6</intersection>
<intersection>195.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>170.5,-478,170.5,-468.5</points>
<intersection>-478 1</intersection>
<intersection>-468.5 8</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>195.5,-478,195.5,-468.5</points>
<intersection>-478 1</intersection>
<intersection>-468.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>170.5,-468.5,196.5,-468.5</points>
<connection>
<GID>231</GID>
<name>clock</name></connection>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<intersection>170.5 6</intersection>
<intersection>195.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179,-476,179.5,-476</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-474,179.5,-470.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>231</GID>
<name>nQ</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-204.5,201,-204.5</points>
<connection>
<GID>224</GID>
<name>N_in0</name></connection>
<connection>
<GID>227</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-465.5,186.5,-462.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<connection>
<GID>235</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-475,186.5,-467.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>-475 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>185.5,-475,186.5,-475</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-470.5,194,-466.5</points>
<intersection>-470.5 3</intersection>
<intersection>-466.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,-466.5,196.5,-466.5</points>
<connection>
<GID>232</GID>
<name>J</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>194,-470.5,196.5,-470.5</points>
<connection>
<GID>232</GID>
<name>K</name></connection>
<intersection>194 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-243.5,185,-209.5</points>
<intersection>-243.5 3</intersection>
<intersection>-209.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-209.5,195,-209.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<connection>
<GID>397</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-243.5,195,-243.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-494,160,-489</points>
<connection>
<GID>253</GID>
<name>clock</name></connection>
<intersection>-494 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-494,160,-494</points>
<intersection>135 2</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>135,-494,135,-484.5</points>
<intersection>-494 1</intersection>
<intersection>-484.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>130.5,-484.5,135,-484.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>135 2</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>159.5,-476.5,159.5,-474</points>
<intersection>-476.5 34</intersection>
<intersection>-474 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>158,-474,161,-474</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>159.5 5</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>159.5,-476.5,160,-476.5</points>
<intersection>159.5 5</intersection>
<intersection>160 41</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>160,-478,160,-476.5</points>
<connection>
<GID>253</GID>
<name>load</name></connection>
<intersection>-476.5 34</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-478,161,-478</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<connection>
<GID>253</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-478,162,-471.5</points>
<connection>
<GID>253</GID>
<name>count_up</name></connection>
<intersection>-471.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-471.5,162,-471.5</points>
<intersection>138 2</intersection>
<intersection>162 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>138,-488.5,138,-468.5</points>
<intersection>-488.5 3</intersection>
<intersection>-471.5 1</intersection>
<intersection>-468.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130.5,-488.5,138,-488.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>138 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>168,-476,168,-461.5</points>
<intersection>-476 6</intersection>
<intersection>-468.5 7</intersection>
<intersection>-461.5 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>168,-476,175,-476</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>168 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>138,-468.5,168,-468.5</points>
<intersection>138 2</intersection>
<intersection>168 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>168,-461.5,180.5,-461.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>168 5</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-520.5,224,-451</points>
<intersection>-520.5 3</intersection>
<intersection>-480 2</intersection>
<intersection>-451 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-451,239,-451</points>
<connection>
<GID>1478</GID>
<name>IN_0</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-480,224,-480</points>
<connection>
<GID>253</GID>
<name>OUT_7</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>224,-520.5,242.5,-520.5</points>
<connection>
<GID>1505</GID>
<name>IN_1</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222,-516.5,222,-447</points>
<intersection>-516.5 3</intersection>
<intersection>-481 2</intersection>
<intersection>-447 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222,-447,239,-447</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-481,222,-481</points>
<connection>
<GID>253</GID>
<name>OUT_6</name></connection>
<intersection>222 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>222,-516.5,242.5,-516.5</points>
<connection>
<GID>1504</GID>
<name>IN_1</name></connection>
<intersection>222 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-512.5,220,-443</points>
<intersection>-512.5 4</intersection>
<intersection>-482 2</intersection>
<intersection>-443 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>220,-443,239,-443</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-482,220,-482</points>
<connection>
<GID>253</GID>
<name>OUT_5</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>220,-512.5,242.5,-512.5</points>
<connection>
<GID>1503</GID>
<name>IN_1</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-508.5,218,-439</points>
<intersection>-508.5 4</intersection>
<intersection>-483 2</intersection>
<intersection>-439 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-439,239,-439</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-483,218,-483</points>
<connection>
<GID>253</GID>
<name>OUT_4</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>218,-508.5,242.5,-508.5</points>
<connection>
<GID>1502</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,-504.5,216,-435</points>
<intersection>-504.5 4</intersection>
<intersection>-484 1</intersection>
<intersection>-435 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-484,216,-484</points>
<connection>
<GID>253</GID>
<name>OUT_3</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-435,239,-435</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>216,-504.5,242.5,-504.5</points>
<connection>
<GID>1501</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-500.5,214,-431</points>
<intersection>-500.5 3</intersection>
<intersection>-485 1</intersection>
<intersection>-431 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-485,214,-485</points>
<connection>
<GID>253</GID>
<name>OUT_2</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-431,239,-431</points>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>214,-500.5,242.5,-500.5</points>
<connection>
<GID>1500</GID>
<name>IN_1</name></connection>
<intersection>214 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-496.5,212,-427</points>
<intersection>-496.5 3</intersection>
<intersection>-486 1</intersection>
<intersection>-427 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-486,212,-486</points>
<connection>
<GID>253</GID>
<name>OUT_1</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212,-427,239,-427</points>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>212,-496.5,242.5,-496.5</points>
<connection>
<GID>1499</GID>
<name>IN_1</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-492.5,210,-423</points>
<intersection>-492.5 3</intersection>
<intersection>-487 1</intersection>
<intersection>-423 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-487,210,-487</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>210,-423,239,-423</points>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>210,-492.5,242.5,-492.5</points>
<connection>
<GID>1498</GID>
<name>IN_1</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306,-450.5,306,-431.5</points>
<intersection>-450.5 1</intersection>
<intersection>-431.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306,-450.5,318,-450.5</points>
<connection>
<GID>1506</GID>
<name>IN_0</name></connection>
<intersection>306 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-431.5,306,-431.5</points>
<connection>
<GID>1426</GID>
<name>N_in1</name></connection>
<intersection>306 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,-449.5,307,-435.5</points>
<intersection>-449.5 1</intersection>
<intersection>-435.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307,-449.5,318,-449.5</points>
<connection>
<GID>1506</GID>
<name>IN_1</name></connection>
<intersection>307 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-435.5,307,-435.5</points>
<connection>
<GID>1428</GID>
<name>N_in1</name></connection>
<intersection>307 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-448.5,308,-439.5</points>
<intersection>-448.5 2</intersection>
<intersection>-439.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-439.5,308,-439.5</points>
<connection>
<GID>1429</GID>
<name>N_in1</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-448.5,318,-448.5</points>
<connection>
<GID>1506</GID>
<name>IN_2</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-447.5,310,-443.5</points>
<intersection>-447.5 2</intersection>
<intersection>-443.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-443.5,310,-443.5</points>
<connection>
<GID>1427</GID>
<name>N_in1</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>310,-447.5,318,-447.5</points>
<connection>
<GID>1506</GID>
<name>IN_3</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-447.5,309,-446.5</points>
<intersection>-447.5 1</intersection>
<intersection>-446.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-447.5,309,-447.5</points>
<connection>
<GID>1430</GID>
<name>N_in1</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-446.5,318,-446.5</points>
<connection>
<GID>1506</GID>
<name>IN_4</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-451.5,313,-445.5</points>
<intersection>-451.5 1</intersection>
<intersection>-445.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-451.5,313,-451.5</points>
<connection>
<GID>1431</GID>
<name>N_in1</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313,-445.5,318,-445.5</points>
<connection>
<GID>1506</GID>
<name>IN_5</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-455.5,312,-444.5</points>
<intersection>-455.5 1</intersection>
<intersection>-444.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-455.5,312,-455.5</points>
<connection>
<GID>1432</GID>
<name>N_in1</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312,-444.5,318,-444.5</points>
<connection>
<GID>1506</GID>
<name>IN_6</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-459.5,311,-443.5</points>
<intersection>-459.5 1</intersection>
<intersection>-443.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-459.5,311,-459.5</points>
<connection>
<GID>1433</GID>
<name>N_in1</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>311,-443.5,318,-443.5</points>
<connection>
<GID>1506</GID>
<name>IN_7</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-482.5,314,-468</points>
<intersection>-482.5 1</intersection>
<intersection>-468 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-482.5,320,-482.5</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-468,314,-468</points>
<connection>
<GID>1434</GID>
<name>N_in1</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-481.5,313,-472</points>
<intersection>-481.5 1</intersection>
<intersection>-472 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-481.5,320,-481.5</points>
<connection>
<GID>1511</GID>
<name>IN_1</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-472,313,-472</points>
<connection>
<GID>1436</GID>
<name>N_in1</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307,-480.5,307,-476</points>
<intersection>-480.5 1</intersection>
<intersection>-476 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>307,-480.5,320,-480.5</points>
<connection>
<GID>1511</GID>
<name>IN_2</name></connection>
<intersection>307 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-476,307,-476</points>
<connection>
<GID>1437</GID>
<name>N_in1</name></connection>
<intersection>307 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-480,311,-479.5</points>
<intersection>-480 2</intersection>
<intersection>-479.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-479.5,320,-479.5</points>
<connection>
<GID>1511</GID>
<name>IN_3</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-480,311,-480</points>
<connection>
<GID>1435</GID>
<name>N_in1</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-484,309,-478.5</points>
<intersection>-484 2</intersection>
<intersection>-478.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-478.5,320,-478.5</points>
<connection>
<GID>1511</GID>
<name>IN_4</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-484,309,-484</points>
<connection>
<GID>1438</GID>
<name>N_in1</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-488,312,-477.5</points>
<intersection>-488 2</intersection>
<intersection>-477.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312,-477.5,320,-477.5</points>
<connection>
<GID>1511</GID>
<name>IN_5</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-488,312,-488</points>
<connection>
<GID>1439</GID>
<name>N_in1</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-492,310,-476.5</points>
<intersection>-492 2</intersection>
<intersection>-476.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-476.5,320,-476.5</points>
<connection>
<GID>1511</GID>
<name>IN_6</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-492,310,-492</points>
<connection>
<GID>1440</GID>
<name>N_in1</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-496,308,-475.5</points>
<intersection>-496 2</intersection>
<intersection>-475.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>308,-475.5,320,-475.5</points>
<connection>
<GID>1511</GID>
<name>IN_7</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,-496,308,-496</points>
<connection>
<GID>1441</GID>
<name>N_in1</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-524,316,-508</points>
<intersection>-524 1</intersection>
<intersection>-508 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-524,322,-524</points>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-508,316,-508</points>
<connection>
<GID>1324</GID>
<name>N_in1</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315,-523,315,-512</points>
<intersection>-523 1</intersection>
<intersection>-512 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315,-523,322,-523</points>
<connection>
<GID>1507</GID>
<name>IN_1</name></connection>
<intersection>315 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-512,315,-512</points>
<connection>
<GID>1326</GID>
<name>N_in1</name></connection>
<intersection>315 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-29.5,191,-29.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-31.5,191,-31.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-33.5,191,-33.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-38,191,-37.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-39.5,191,-39.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-41.5,191,-41.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-43.5,191,-43.5</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-35.5,191,-35.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-522,310,-516</points>
<intersection>-522 1</intersection>
<intersection>-516 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-522,322,-522</points>
<connection>
<GID>1507</GID>
<name>IN_2</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-516,310,-516</points>
<connection>
<GID>1327</GID>
<name>N_in1</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-521,309,-520</points>
<intersection>-521 1</intersection>
<intersection>-520 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-521,322,-521</points>
<connection>
<GID>1507</GID>
<name>IN_3</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-520,309,-520</points>
<connection>
<GID>1325</GID>
<name>N_in1</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313,-524,313,-520</points>
<intersection>-524 2</intersection>
<intersection>-520 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313,-520,322,-520</points>
<connection>
<GID>1507</GID>
<name>IN_4</name></connection>
<intersection>313 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-524,313,-524</points>
<connection>
<GID>1328</GID>
<name>N_in1</name></connection>
<intersection>313 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312,-528,312,-519</points>
<intersection>-528 2</intersection>
<intersection>-519 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312,-519,322,-519</points>
<connection>
<GID>1507</GID>
<name>IN_5</name></connection>
<intersection>312 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-528,312,-528</points>
<connection>
<GID>1329</GID>
<name>N_in1</name></connection>
<intersection>312 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-532,314,-518</points>
<intersection>-532 2</intersection>
<intersection>-518 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-518,322,-518</points>
<connection>
<GID>1507</GID>
<name>IN_6</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-532,314,-532</points>
<connection>
<GID>1330</GID>
<name>N_in1</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-536,311,-517</points>
<intersection>-536 2</intersection>
<intersection>-517 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-517,322,-517</points>
<connection>
<GID>1507</GID>
<name>IN_7</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,-536,311,-536</points>
<connection>
<GID>1331</GID>
<name>N_in1</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-247.5,185.5,-213.5</points>
<intersection>-247.5 3</intersection>
<intersection>-213.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>176,-213.5,195,-213.5</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>398</GID>
<name>OUT</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185.5,-247.5,195,-247.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>186,-251.5,186,-217.5</points>
<intersection>-251.5 5</intersection>
<intersection>-217.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>186,-251.5,195,-251.5</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<intersection>186 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>176,-217.5,195,-217.5</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<intersection>186 4</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>186.5,-255.5,186.5,-221.5</points>
<intersection>-255.5 4</intersection>
<intersection>-221.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>186.5,-255.5,195,-255.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>186.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>176,-221.5,195,-221.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>186.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>187.5,-225.5,195,-225.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>187.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>187.5,-259.5,187.5,-225.5</points>
<intersection>-259.5 4</intersection>
<intersection>-226.5 5</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>187.5,-259.5,195,-259.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>187.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>170,-226.5,187.5,-226.5</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<intersection>187.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>176,-229.5,195,-229.5</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<intersection>187.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>187.5,-263.5,187.5,-229.5</points>
<intersection>-263.5 4</intersection>
<intersection>-229.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>187.5,-263.5,195,-263.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>187.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>188,-267.5,188,-233.5</points>
<intersection>-267.5 4</intersection>
<intersection>-233.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>188,-267.5,195,-267.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>188 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>176,-233.5,195,-233.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>188 3</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-212.5,201,-212.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-208.5,201,-208.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<connection>
<GID>257</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-216.5,201,-216.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<connection>
<GID>255</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-220.5,201,-220.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<connection>
<GID>259</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-224.5,201,-224.5</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<connection>
<GID>260</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-228.5,201,-228.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<connection>
<GID>261</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-232.5,201,-232.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<connection>
<GID>270</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>201,-238.5,201,-238.5</points>
<connection>
<GID>271</GID>
<name>N_in0</name></connection>
<connection>
<GID>272</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-246.5,201,-246.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<connection>
<GID>282</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-242.5,201,-242.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<connection>
<GID>281</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-250.5,201,-250.5</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<connection>
<GID>280</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-254.5,201,-254.5</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<connection>
<GID>283</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-258.5,201,-258.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<connection>
<GID>284</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-262.5,201,-262.5</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>285</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-266.5,201,-266.5</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>286</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-231.5,195,-231.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-227.5,195,-227.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<connection>
<GID>292</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-223.5,195,-223.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-219.5,195,-219.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-215.5,195,-215.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-211.5,195,-211.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-207.5,195,-207.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-273,195,-273</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>184.5,-309,184.5,-275</points>
<intersection>-309 19</intersection>
<intersection>-275 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>175.5,-275,195,-275</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<connection>
<GID>415</GID>
<name>OUT</name></connection>
<intersection>184.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>184.5,-309,195,-309</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>184.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>201,-274,201,-274</points>
<connection>
<GID>295</GID>
<name>N_in0</name></connection>
<connection>
<GID>296</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-313,185,-279</points>
<intersection>-313 3</intersection>
<intersection>-279 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-279,195,-279</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185,-313,195,-313</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-317,185.5,-283</points>
<intersection>-317 3</intersection>
<intersection>-283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-283,195,-283</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185.5,-317,195,-317</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>186,-321,186,-287</points>
<intersection>-321 5</intersection>
<intersection>-287 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>186,-321,195,-321</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>186 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>175.5,-287,195,-287</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>186 4</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>186.5,-325,186.5,-291</points>
<intersection>-325 4</intersection>
<intersection>-291 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>186.5,-325,195,-325</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>186.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>175.5,-291,195,-291</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<connection>
<GID>419</GID>
<name>OUT</name></connection>
<intersection>186.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>187,-329,187,-295</points>
<intersection>-329 4</intersection>
<intersection>-295 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>187,-329,195,-329</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>187 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>175.5,-295,195,-295</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<connection>
<GID>420</GID>
<name>OUT</name></connection>
<intersection>187 3</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175.5,-299,195,-299</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<intersection>187.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>187.5,-333,187.5,-299</points>
<intersection>-333 4</intersection>
<intersection>-299 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>187.5,-333,195,-333</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>187.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>188,-337,188,-303</points>
<intersection>-337 4</intersection>
<intersection>-303 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>188,-337,195,-337</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>188 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>175.5,-303,195,-303</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<connection>
<GID>422</GID>
<name>OUT</name></connection>
<intersection>188 3</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-282,201,-282</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<connection>
<GID>307</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-278,201,-278</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-286,201,-286</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<connection>
<GID>305</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-290,201,-290</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<connection>
<GID>308</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-294,201,-294</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>309</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-298,201,-298</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<connection>
<GID>310</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-302,201,-302</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<connection>
<GID>311</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>201,-308,201,-308</points>
<connection>
<GID>312</GID>
<name>N_in0</name></connection>
<connection>
<GID>313</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-316,201,-316</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<connection>
<GID>323</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-312,201,-312</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<connection>
<GID>322</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-320,201,-320</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<connection>
<GID>321</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-324,201,-324</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<connection>
<GID>325</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-328,201,-328</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<connection>
<GID>327</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-332,201,-332</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<connection>
<GID>329</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-336,201,-336</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<connection>
<GID>332</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-301,195,-301</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-335,184,-197.5</points>
<intersection>-335 18</intersection>
<intersection>-331 17</intersection>
<intersection>-327 16</intersection>
<intersection>-323 15</intersection>
<intersection>-319 14</intersection>
<intersection>-315 13</intersection>
<intersection>-311 12</intersection>
<intersection>-307 11</intersection>
<intersection>-301 2</intersection>
<intersection>-297 9</intersection>
<intersection>-293 8</intersection>
<intersection>-289 7</intersection>
<intersection>-285 6</intersection>
<intersection>-281 5</intersection>
<intersection>-277 4</intersection>
<intersection>-273 3</intersection>
<intersection>-265.5 38</intersection>
<intersection>-261.5 37</intersection>
<intersection>-257.5 36</intersection>
<intersection>-253.5 35</intersection>
<intersection>-249.5 34</intersection>
<intersection>-245.5 33</intersection>
<intersection>-241.5 32</intersection>
<intersection>-237.5 31</intersection>
<intersection>-231.5 22</intersection>
<intersection>-227.5 29</intersection>
<intersection>-223.5 28</intersection>
<intersection>-219.5 27</intersection>
<intersection>-215.5 26</intersection>
<intersection>-211.5 25</intersection>
<intersection>-207.5 24</intersection>
<intersection>-203.5 23</intersection>
<intersection>-197.5 21</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>184,-301,191,-301</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184,-273,191,-273</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>184,-277,191,-277</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>184,-281,191,-281</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>184,-285,191,-285</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>184,-289,191,-289</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>184,-293,191,-293</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>184,-297,191,-297</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>184,-307,195,-307</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>184,-311,195,-311</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>184,-315,195,-315</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>184,-319,195,-319</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>184,-323,195,-323</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>184,-327,195,-327</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>184,-331,195,-331</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>184,-335,195,-335</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>146.5,-197.5,184,-197.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>184,-231.5,191,-231.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>184,-203.5,191,-203.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>184,-207.5,191,-207.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>184,-211.5,191,-211.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>184,-215.5,191,-215.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>184,-219.5,191,-219.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>184,-223.5,191,-223.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>184,-227.5,191,-227.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>184,-237.5,195,-237.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>184,-241.5,195,-241.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>184,-245.5,195,-245.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>184,-249.5,195,-249.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>184,-253.5,195,-253.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>184,-257.5,195,-257.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>184,-261.5,195,-261.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>184,-265.5,195,-265.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-297,195,-297</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-293,195,-293</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-289,195,-289</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-285,195,-285</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-281,195,-281</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>195,-277,195,-277</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-251.5,229,-251.5</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>348</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-255.5,229,-255.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<connection>
<GID>350</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-279.5,229,-279.5</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<connection>
<GID>355</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-259.5,229,-259.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>351</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-263.5,229,-263.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>349</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-267.5,229,-267.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>352</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-271.5,229,-271.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>353</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-275.5,229,-275.5</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<connection>
<GID>354</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-215,227,-204.5</points>
<intersection>-215 1</intersection>
<intersection>-204.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-215,229,-215</points>
<connection>
<GID>340</GID>
<name>N_in0</name></connection>
<intersection>227 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-204.5,227,-204.5</points>
<connection>
<GID>224</GID>
<name>N_in1</name></connection>
<intersection>227 0</intersection></hsegment></shape></wire>
<wire>
<ID>1021</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-240,42,-239.5</points>
<connection>
<GID>1259</GID>
<name>IN_0</name></connection>
<connection>
<GID>1256</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-219,225.5,-208.5</points>
<intersection>-219 2</intersection>
<intersection>-208.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-208.5,225.5,-208.5</points>
<connection>
<GID>257</GID>
<name>N_in1</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-219,229,-219</points>
<connection>
<GID>342</GID>
<name>N_in0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1022</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-243.5,42,-243.5</points>
<connection>
<GID>1260</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-223,224,-212.5</points>
<intersection>-223 2</intersection>
<intersection>-212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-212.5,224,-212.5</points>
<connection>
<GID>258</GID>
<name>N_in1</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>224,-223,229,-223</points>
<connection>
<GID>343</GID>
<name>N_in0</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-245.5,42,-245.5</points>
<connection>
<GID>1262</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-227,222.5,-216.5</points>
<intersection>-227 1</intersection>
<intersection>-216.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-227,229,-227</points>
<connection>
<GID>341</GID>
<name>N_in0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-216.5,222.5,-216.5</points>
<connection>
<GID>255</GID>
<name>N_in1</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-247.5,42,-247.5</points>
<connection>
<GID>1264</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,-231,221.5,-220.5</points>
<intersection>-231 1</intersection>
<intersection>-220.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221.5,-231,229,-231</points>
<connection>
<GID>344</GID>
<name>N_in0</name></connection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-220.5,221.5,-220.5</points>
<connection>
<GID>259</GID>
<name>N_in1</name></connection>
<intersection>221.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1025</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>42,-249.5,42,-249.5</points>
<connection>
<GID>1266</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-235,220,-224.5</points>
<intersection>-235 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-224.5,220,-224.5</points>
<connection>
<GID>260</GID>
<name>N_in1</name></connection>
<intersection>220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-235,229,-235</points>
<connection>
<GID>345</GID>
<name>N_in0</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>1026</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-251.5,42,-251.5</points>
<connection>
<GID>1268</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1269</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-239,219,-228.5</points>
<intersection>-239 1</intersection>
<intersection>-228.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-239,229,-239</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-228.5,219,-228.5</points>
<connection>
<GID>261</GID>
<name>N_in1</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>1027</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-253.5,42,-253.5</points>
<connection>
<GID>1270</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-243,218,-232.5</points>
<intersection>-243 2</intersection>
<intersection>-232.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-232.5,218,-232.5</points>
<connection>
<GID>270</GID>
<name>N_in1</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,-243,229,-243</points>
<connection>
<GID>347</GID>
<name>N_in0</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>1028</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-255.5,42,-255.5</points>
<connection>
<GID>1272</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1273</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,-250.5,216,-238.5</points>
<intersection>-250.5 1</intersection>
<intersection>-238.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,-250.5,223,-250.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-238.5,216,-238.5</points>
<connection>
<GID>271</GID>
<name>N_in1</name></connection>
<intersection>216 0</intersection></hsegment></shape></wire>
<wire>
<ID>1029</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-257.5,42,-257.5</points>
<connection>
<GID>1274</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1275</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-254.5,214.5,-242.5</points>
<intersection>-254.5 1</intersection>
<intersection>-242.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>214.5,-254.5,223,-254.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>214.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-242.5,214.5,-242.5</points>
<connection>
<GID>281</GID>
<name>N_in1</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1030</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-203,70.5,-203</points>
<connection>
<GID>1276</GID>
<name>IN_0</name></connection>
<connection>
<GID>1278</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-258.5,213,-246.5</points>
<intersection>-258.5 1</intersection>
<intersection>-246.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-258.5,223,-258.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-246.5,213,-246.5</points>
<connection>
<GID>282</GID>
<name>N_in1</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>1031</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-207,70.5,-207</points>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection>
<connection>
<GID>1280</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-262.5,211.5,-250.5</points>
<intersection>-262.5 1</intersection>
<intersection>-250.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-262.5,223,-262.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-250.5,211.5,-250.5</points>
<connection>
<GID>280</GID>
<name>N_in1</name></connection>
<intersection>211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1032</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-211,70.5,-211</points>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection>
<connection>
<GID>1282</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-266.5,210,-254.5</points>
<intersection>-266.5 1</intersection>
<intersection>-254.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210,-266.5,223,-266.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-254.5,210,-254.5</points>
<connection>
<GID>283</GID>
<name>N_in1</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>1033</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-215,70.5,-215</points>
<connection>
<GID>1283</GID>
<name>IN_0</name></connection>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,-270.5,208.5,-258.5</points>
<intersection>-270.5 1</intersection>
<intersection>-258.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-270.5,223,-270.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-258.5,208.5,-258.5</points>
<connection>
<GID>284</GID>
<name>N_in1</name></connection>
<intersection>208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1034</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-219,70.5,-219</points>
<connection>
<GID>1285</GID>
<name>IN_0</name></connection>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-274.5,207,-262.5</points>
<intersection>-274.5 1</intersection>
<intersection>-262.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-274.5,223,-274.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-262.5,207,-262.5</points>
<connection>
<GID>285</GID>
<name>N_in1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>1035</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-223,70.5,-223</points>
<connection>
<GID>1287</GID>
<name>IN_0</name></connection>
<connection>
<GID>1288</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-278.5,205.5,-266.5</points>
<intersection>-278.5 1</intersection>
<intersection>-266.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-278.5,223,-278.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>205.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-266.5,205.5,-266.5</points>
<connection>
<GID>286</GID>
<name>N_in1</name></connection>
<intersection>205.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1036</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-227,70.5,-227</points>
<connection>
<GID>1289</GID>
<name>IN_0</name></connection>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-274,217,-252.5</points>
<intersection>-274 2</intersection>
<intersection>-252.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-252.5,223,-252.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-274,217,-274</points>
<connection>
<GID>295</GID>
<name>N_in1</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>1037</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-231,70.5,-231</points>
<connection>
<GID>1291</GID>
<name>IN_0</name></connection>
<connection>
<GID>1292</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-278,215.5,-256.5</points>
<intersection>-278 1</intersection>
<intersection>-256.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-278,215.5,-278</points>
<connection>
<GID>306</GID>
<name>N_in1</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>215.5,-256.5,223,-256.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1038</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-203,74.5,-203</points>
<connection>
<GID>1278</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1293</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214,-282,214,-260.5</points>
<intersection>-282 1</intersection>
<intersection>-260.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-282,214,-282</points>
<connection>
<GID>307</GID>
<name>N_in1</name></connection>
<intersection>214 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-260.5,223,-260.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>214 0</intersection></hsegment></shape></wire>
<wire>
<ID>1039</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-207,74.5,-207</points>
<connection>
<GID>1280</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1294</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,-286,212.5,-264.5</points>
<intersection>-286 1</intersection>
<intersection>-264.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-286,212.5,-286</points>
<connection>
<GID>305</GID>
<name>N_in1</name></connection>
<intersection>212.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>212.5,-264.5,223,-264.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>212.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1040</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-211,74.5,-211</points>
<connection>
<GID>1282</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1295</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-290,211,-268.5</points>
<intersection>-290 1</intersection>
<intersection>-268.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-290,211,-290</points>
<connection>
<GID>308</GID>
<name>N_in1</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>211,-268.5,223,-268.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>1041</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-215,74.5,-215</points>
<connection>
<GID>1284</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1296</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209.5,-294,209.5,-272.5</points>
<intersection>-294 1</intersection>
<intersection>-272.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-294,209.5,-294</points>
<connection>
<GID>309</GID>
<name>N_in1</name></connection>
<intersection>209.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209.5,-272.5,223,-272.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>209.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1042</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-219,74.5,-219</points>
<connection>
<GID>1286</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1297</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-298,208,-276.5</points>
<intersection>-298 1</intersection>
<intersection>-276.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-298,208,-298</points>
<connection>
<GID>310</GID>
<name>N_in1</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>208,-276.5,223,-276.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>1043</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-223,74.5,-223</points>
<connection>
<GID>1288</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1298</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206.5,-302,206.5,-280.5</points>
<intersection>-302 1</intersection>
<intersection>-280.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-302,206.5,-302</points>
<connection>
<GID>311</GID>
<name>N_in1</name></connection>
<intersection>206.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206.5,-280.5,223,-280.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>206.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1044</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-227,74.5,-227</points>
<connection>
<GID>1290</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1299</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-308,213.5,-291.5</points>
<intersection>-308 2</intersection>
<intersection>-291.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-291.5,229.5,-291.5</points>
<connection>
<GID>4</GID>
<name>N_in0</name></connection>
<intersection>213.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-308,213.5,-308</points>
<connection>
<GID>312</GID>
<name>N_in1</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1045</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-231,74.5,-231</points>
<connection>
<GID>1292</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1300</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-312,215.5,-295.5</points>
<intersection>-312 2</intersection>
<intersection>-295.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-295.5,229.5,-295.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<intersection>215.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-312,215.5,-312</points>
<connection>
<GID>322</GID>
<name>N_in1</name></connection>
<intersection>215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1046</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-201,58.5,-201</points>
<connection>
<GID>1258</GID>
<name>IN_0</name></connection>
<connection>
<GID>1301</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217,-316,217,-299.5</points>
<intersection>-316 2</intersection>
<intersection>-299.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217,-299.5,229.5,-299.5</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>217 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-316,217,-316</points>
<connection>
<GID>323</GID>
<name>N_in1</name></connection>
<intersection>217 0</intersection></hsegment></shape></wire>
<wire>
<ID>1047</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-201,74.5,-201</points>
<connection>
<GID>1293</GID>
<name>IN_0</name></connection>
<connection>
<GID>1301</GID>
<name>OUT_0</name></connection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-229,63,-201</points>
<intersection>-229 4</intersection>
<intersection>-225 10</intersection>
<intersection>-221 9</intersection>
<intersection>-217 8</intersection>
<intersection>-213 7</intersection>
<intersection>-209 6</intersection>
<intersection>-205 5</intersection>
<intersection>-201 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63,-229,74.5,-229</points>
<connection>
<GID>1300</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-205,74.5,-205</points>
<connection>
<GID>1294</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63,-209,74.5,-209</points>
<connection>
<GID>1295</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>63,-213,74.5,-213</points>
<connection>
<GID>1296</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>63,-217,74.5,-217</points>
<connection>
<GID>1297</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>63,-221,74.5,-221</points>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>63,-225,74.5,-225</points>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection>
<intersection>63 3</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-320,219,-303.5</points>
<intersection>-320 2</intersection>
<intersection>-303.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-303.5,229.5,-303.5</points>
<connection>
<GID>15</GID>
<name>N_in0</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-320,219,-320</points>
<connection>
<GID>321</GID>
<name>N_in1</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>1048</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-237,74.5,-237</points>
<connection>
<GID>1302</GID>
<name>IN_0</name></connection>
<connection>
<GID>1312</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68.5,-265,68.5,-237</points>
<intersection>-265 4</intersection>
<intersection>-261 10</intersection>
<intersection>-257 9</intersection>
<intersection>-253 8</intersection>
<intersection>-249 7</intersection>
<intersection>-245 6</intersection>
<intersection>-241 5</intersection>
<intersection>-237 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-265,74.5,-265</points>
<connection>
<GID>1319</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-241,74.5,-241</points>
<connection>
<GID>1313</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>68.5,-245,74.5,-245</points>
<connection>
<GID>1314</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,-249,74.5,-249</points>
<connection>
<GID>1315</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>68.5,-253,74.5,-253</points>
<connection>
<GID>1316</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>68.5,-257,74.5,-257</points>
<connection>
<GID>1317</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>68.5,-261,74.5,-261</points>
<connection>
<GID>1318</GID>
<name>IN_0</name></connection>
<intersection>68.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221,-324,221,-307.5</points>
<intersection>-324 2</intersection>
<intersection>-307.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221,-307.5,229.5,-307.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>221 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-324,221,-324</points>
<connection>
<GID>325</GID>
<name>N_in1</name></connection>
<intersection>221 0</intersection></hsegment></shape></wire>
<wire>
<ID>1049</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-239,74.5,-239</points>
<connection>
<GID>1303</GID>
<name>IN_0</name></connection>
<connection>
<GID>1312</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,-328,223.5,-311.5</points>
<intersection>-328 2</intersection>
<intersection>-311.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,-311.5,229.5,-311.5</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<intersection>223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-328,223.5,-328</points>
<connection>
<GID>327</GID>
<name>N_in1</name></connection>
<intersection>223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1050</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-243,74.5,-243</points>
<connection>
<GID>1305</GID>
<name>IN_0</name></connection>
<connection>
<GID>1313</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-332,225.5,-315.5</points>
<intersection>-332 1</intersection>
<intersection>-315.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>203,-332,225.5,-332</points>
<connection>
<GID>329</GID>
<name>N_in1</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-315.5,229.5,-315.5</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1051</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-247,74.5,-247</points>
<connection>
<GID>1306</GID>
<name>IN_0</name></connection>
<connection>
<GID>1314</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,-336,227.5,-319.5</points>
<intersection>-336 2</intersection>
<intersection>-319.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,-319.5,229.5,-319.5</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203,-336,227.5,-336</points>
<connection>
<GID>332</GID>
<name>N_in1</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1052</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-251,74.5,-251</points>
<connection>
<GID>1307</GID>
<name>IN_0</name></connection>
<connection>
<GID>1315</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1053</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-255,74.5,-255</points>
<connection>
<GID>1308</GID>
<name>IN_0</name></connection>
<connection>
<GID>1316</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1054</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-267,74.5,-267</points>
<connection>
<GID>1311</GID>
<name>IN_0</name></connection>
<connection>
<GID>1319</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1055</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-263,74.5,-263</points>
<connection>
<GID>1310</GID>
<name>IN_0</name></connection>
<connection>
<GID>1318</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1056</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-259,74.5,-259</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<connection>
<GID>1317</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1061</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-420,268,-420</points>
<connection>
<GID>1346</GID>
<name>IN_0</name></connection>
<connection>
<GID>1347</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-206.5,166,-206.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1062</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>257.5,-456,257.5,-422</points>
<intersection>-456 19</intersection>
<intersection>-422 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>249,-422,268,-422</points>
<connection>
<GID>1346</GID>
<name>IN_1</name></connection>
<connection>
<GID>1479</GID>
<name>OUT</name></connection>
<intersection>257.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>257.5,-456,268,-456</points>
<connection>
<GID>1363</GID>
<name>IN_1</name></connection>
<intersection>257.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-210.5,166,-210.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<connection>
<GID>380</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1063</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-421,274,-421</points>
<connection>
<GID>1345</GID>
<name>N_in0</name></connection>
<connection>
<GID>1346</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-214.5,166,-214.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1064</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-460,258,-426</points>
<intersection>-460 3</intersection>
<intersection>-426 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249,-426,268,-426</points>
<connection>
<GID>1348</GID>
<name>IN_1</name></connection>
<connection>
<GID>1480</GID>
<name>OUT</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258,-460,268,-460</points>
<connection>
<GID>1364</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-218.5,166,-218.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1065</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-464,258.5,-430</points>
<intersection>-464 3</intersection>
<intersection>-430 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249,-430,268,-430</points>
<connection>
<GID>1349</GID>
<name>IN_1</name></connection>
<connection>
<GID>1481</GID>
<name>OUT</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,-464,268,-464</points>
<connection>
<GID>1365</GID>
<name>IN_1</name></connection>
<intersection>258.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-222.5,166,-222.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1066</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>259,-468,259,-434</points>
<intersection>-468 5</intersection>
<intersection>-434 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>259,-468,268,-468</points>
<connection>
<GID>1366</GID>
<name>IN_1</name></connection>
<intersection>259 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>249,-434,268,-434</points>
<connection>
<GID>1350</GID>
<name>IN_1</name></connection>
<connection>
<GID>1482</GID>
<name>OUT</name></connection>
<intersection>259 4</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-226.5,166,-226.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1067</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>259.5,-472,259.5,-438</points>
<intersection>-472 4</intersection>
<intersection>-438 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-472,268,-472</points>
<connection>
<GID>1367</GID>
<name>IN_1</name></connection>
<intersection>259.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>249,-438,268,-438</points>
<connection>
<GID>1351</GID>
<name>IN_1</name></connection>
<connection>
<GID>1483</GID>
<name>OUT</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-230.5,166,-230.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1068</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>249,-442,268,-442</points>
<connection>
<GID>1352</GID>
<name>IN_1</name></connection>
<connection>
<GID>1484</GID>
<name>OUT</name></connection>
<intersection>258 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>258,-476,258,-442</points>
<intersection>-476 4</intersection>
<intersection>-442 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258,-476,268,-476</points>
<connection>
<GID>1368</GID>
<name>IN_1</name></connection>
<intersection>258 3</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-234.5,166,-234.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1069</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>249,-446,268,-446</points>
<connection>
<GID>1353</GID>
<name>IN_1</name></connection>
<connection>
<GID>1485</GID>
<name>OUT</name></connection>
<intersection>258.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>258.5,-480,258.5,-446</points>
<intersection>-480 4</intersection>
<intersection>-446 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258.5,-480,268,-480</points>
<connection>
<GID>1369</GID>
<name>IN_1</name></connection>
<intersection>258.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-206.5,170,-206.5</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<connection>
<GID>395</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1070</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>261,-484,261,-450</points>
<intersection>-484 4</intersection>
<intersection>-450 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,-484,268,-484</points>
<connection>
<GID>1370</GID>
<name>IN_1</name></connection>
<intersection>261 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>249,-450,268,-450</points>
<connection>
<GID>1354</GID>
<name>IN_1</name></connection>
<connection>
<GID>1486</GID>
<name>OUT</name></connection>
<intersection>261 3</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-210.5,170,-210.5</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<connection>
<GID>397</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1071</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-429,274,-429</points>
<connection>
<GID>1349</GID>
<name>OUT</name></connection>
<connection>
<GID>1357</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-214.5,170,-214.5</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<connection>
<GID>398</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1072</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-425,274,-425</points>
<connection>
<GID>1348</GID>
<name>OUT</name></connection>
<connection>
<GID>1356</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-218.5,170,-218.5</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<connection>
<GID>399</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1073</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-433,274,-433</points>
<connection>
<GID>1350</GID>
<name>OUT</name></connection>
<connection>
<GID>1355</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-222.5,170,-222.5</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<connection>
<GID>400</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1074</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-437,274,-437</points>
<connection>
<GID>1351</GID>
<name>OUT</name></connection>
<connection>
<GID>1358</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-230.5,170,-230.5</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1075</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-441,274,-441</points>
<connection>
<GID>1352</GID>
<name>OUT</name></connection>
<connection>
<GID>1359</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-234.5,170,-234.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<connection>
<GID>402</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1076</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-445,274,-445</points>
<connection>
<GID>1353</GID>
<name>OUT</name></connection>
<connection>
<GID>1360</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-204.5,154,-204.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1077</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-449,274,-449</points>
<connection>
<GID>1354</GID>
<name>OUT</name></connection>
<connection>
<GID>1361</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>158,-204.5,170,-204.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>OUT_0</name></connection>
<intersection>158 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158,-232.5,158,-204.5</points>
<intersection>-232.5 4</intersection>
<intersection>-228.5 10</intersection>
<intersection>-220.5 8</intersection>
<intersection>-216.5 7</intersection>
<intersection>-212.5 6</intersection>
<intersection>-208.5 5</intersection>
<intersection>-204.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>158,-232.5,170,-232.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>158,-208.5,170,-208.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>158,-212.5,170,-212.5</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>158,-216.5,170,-216.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>158,-220.5,170,-220.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>158,-228.5,170,-228.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>158 3</intersection></hsegment></shape></wire>
<wire>
<ID>1078</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>274,-455,274,-455</points>
<connection>
<GID>1362</GID>
<name>N_in0</name></connection>
<connection>
<GID>1363</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163.5,-274,169.5,-274</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>163.5,-302,163.5,-274</points>
<intersection>-302 4</intersection>
<intersection>-298 10</intersection>
<intersection>-294 9</intersection>
<intersection>-290 8</intersection>
<intersection>-286 7</intersection>
<intersection>-282 6</intersection>
<intersection>-278 5</intersection>
<intersection>-274 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>163.5,-302,169.5,-302</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>163.5,-278,169.5,-278</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>163.5,-282,169.5,-282</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>163.5,-286,169.5,-286</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>163.5,-290,169.5,-290</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>163.5,-294,169.5,-294</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>163.5,-298,169.5,-298</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>163.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1079</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-463,274,-463</points>
<connection>
<GID>1365</GID>
<name>OUT</name></connection>
<connection>
<GID>1373</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-276,169.5,-276</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<connection>
<GID>415</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1080</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-459,274,-459</points>
<connection>
<GID>1364</GID>
<name>OUT</name></connection>
<connection>
<GID>1372</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1081</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-467,274,-467</points>
<connection>
<GID>1366</GID>
<name>OUT</name></connection>
<connection>
<GID>1371</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,52.5,73.5,72</points>
<intersection>52.5 8</intersection>
<intersection>58.5 1</intersection>
<intersection>72 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,58.5,73.5,58.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>73.5,72,110,72</points>
<connection>
<GID>1515</GID>
<name>clock</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>73.5,52.5,98.5,52.5</points>
<intersection>73.5 0</intersection>
<intersection>98.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>98.5,52.5,98.5,54</points>
<connection>
<GID>1521</GID>
<name>clock</name></connection>
<intersection>52.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-280,169.5,-280</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1082</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-471,274,-471</points>
<connection>
<GID>1367</GID>
<name>OUT</name></connection>
<connection>
<GID>1374</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-284,169.5,-284</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<connection>
<GID>417</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1083</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-475,274,-475</points>
<connection>
<GID>1368</GID>
<name>OUT</name></connection>
<connection>
<GID>1375</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-288,169.5,-288</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<connection>
<GID>418</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1084</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-479,274,-479</points>
<connection>
<GID>1369</GID>
<name>OUT</name></connection>
<connection>
<GID>1376</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-292,169.5,-292</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<connection>
<GID>419</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1085</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-483,274,-483</points>
<connection>
<GID>1370</GID>
<name>OUT</name></connection>
<connection>
<GID>1377</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-304,169.5,-304</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<connection>
<GID>422</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1086</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-448,268,-448</points>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection>
<connection>
<GID>1384</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-300,169.5,-300</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<connection>
<GID>421</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1087</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-444,268,-444</points>
<connection>
<GID>1353</GID>
<name>IN_0</name></connection>
<connection>
<GID>1383</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-296,169.5,-296</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<connection>
<GID>420</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1088</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-440,268,-440</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<connection>
<GID>1382</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1089</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-436,268,-436</points>
<connection>
<GID>1351</GID>
<name>IN_0</name></connection>
<connection>
<GID>1381</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1090</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-432,268,-432</points>
<connection>
<GID>1350</GID>
<name>IN_0</name></connection>
<connection>
<GID>1380</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>98,65,98,69</points>
<intersection>65 34</intersection>
<intersection>69 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>96.5,69,99.5,69</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<connection>
<GID>1519</GID>
<name>OUT_0</name></connection>
<intersection>98 5</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>98,65,98.5,65</points>
<connection>
<GID>1521</GID>
<name>load</name></connection>
<intersection>98 5</intersection></hsegment></shape></wire>
<wire>
<ID>1091</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-428,268,-428</points>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection>
<connection>
<GID>1379</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1092</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-424,268,-424</points>
<connection>
<GID>1348</GID>
<name>IN_0</name></connection>
<connection>
<GID>1378</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1093</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-489.5,268,-489.5</points>
<connection>
<GID>1387</GID>
<name>IN_0</name></connection>
<connection>
<GID>1388</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1094</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>257.5,-525.5,257.5,-491.5</points>
<intersection>-525.5 19</intersection>
<intersection>-491.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>248.5,-491.5,268,-491.5</points>
<connection>
<GID>1387</GID>
<name>IN_1</name></connection>
<connection>
<GID>1498</GID>
<name>OUT</name></connection>
<intersection>257.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>257.5,-525.5,268,-525.5</points>
<connection>
<GID>1404</GID>
<name>IN_1</name></connection>
<intersection>257.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1095</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>274,-490.5,274,-490.5</points>
<connection>
<GID>1386</GID>
<name>N_in0</name></connection>
<connection>
<GID>1387</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1096</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-529.5,258,-495.5</points>
<intersection>-529.5 3</intersection>
<intersection>-495.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248.5,-495.5,268,-495.5</points>
<connection>
<GID>1389</GID>
<name>IN_1</name></connection>
<connection>
<GID>1499</GID>
<name>OUT</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258,-529.5,268,-529.5</points>
<connection>
<GID>1405</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>1097</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-533.5,258.5,-499.5</points>
<intersection>-533.5 3</intersection>
<intersection>-499.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248.5,-499.5,268,-499.5</points>
<connection>
<GID>1390</GID>
<name>IN_1</name></connection>
<connection>
<GID>1500</GID>
<name>OUT</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>258.5,-533.5,268,-533.5</points>
<connection>
<GID>1406</GID>
<name>IN_1</name></connection>
<intersection>258.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1098</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>259,-537.5,259,-503.5</points>
<intersection>-537.5 5</intersection>
<intersection>-503.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>259,-537.5,268,-537.5</points>
<connection>
<GID>1407</GID>
<name>IN_1</name></connection>
<intersection>259 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>248.5,-503.5,268,-503.5</points>
<connection>
<GID>1391</GID>
<name>IN_1</name></connection>
<connection>
<GID>1501</GID>
<name>OUT</name></connection>
<intersection>259 4</intersection></hsegment></shape></wire>
<wire>
<ID>1099</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>259.5,-541.5,259.5,-507.5</points>
<intersection>-541.5 4</intersection>
<intersection>-507.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>259.5,-541.5,268,-541.5</points>
<connection>
<GID>1408</GID>
<name>IN_1</name></connection>
<intersection>259.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>248.5,-507.5,268,-507.5</points>
<connection>
<GID>1392</GID>
<name>IN_1</name></connection>
<connection>
<GID>1502</GID>
<name>OUT</name></connection>
<intersection>259.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1100</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>260,-545.5,260,-511.5</points>
<intersection>-545.5 4</intersection>
<intersection>-511.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>260,-545.5,268,-545.5</points>
<connection>
<GID>1409</GID>
<name>IN_1</name></connection>
<intersection>260 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>248.5,-511.5,268,-511.5</points>
<connection>
<GID>1393</GID>
<name>IN_1</name></connection>
<connection>
<GID>1503</GID>
<name>OUT</name></connection>
<intersection>260 3</intersection></hsegment></shape></wire>
<wire>
<ID>1101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>248.5,-515.5,268,-515.5</points>
<connection>
<GID>1394</GID>
<name>IN_1</name></connection>
<connection>
<GID>1504</GID>
<name>OUT</name></connection>
<intersection>258.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>258.5,-549.5,258.5,-515.5</points>
<intersection>-549.5 4</intersection>
<intersection>-515.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>258.5,-549.5,268,-549.5</points>
<connection>
<GID>1410</GID>
<name>IN_1</name></connection>
<intersection>258.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1102</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>261,-553.5,261,-519.5</points>
<intersection>-553.5 4</intersection>
<intersection>-519.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>261,-553.5,268,-553.5</points>
<connection>
<GID>1411</GID>
<name>IN_1</name></connection>
<intersection>261 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>248.5,-519.5,268,-519.5</points>
<connection>
<GID>1395</GID>
<name>IN_1</name></connection>
<connection>
<GID>1505</GID>
<name>OUT</name></connection>
<intersection>261 3</intersection></hsegment></shape></wire>
<wire>
<ID>1103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-498.5,274,-498.5</points>
<connection>
<GID>1390</GID>
<name>OUT</name></connection>
<connection>
<GID>1398</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-494.5,274,-494.5</points>
<connection>
<GID>1389</GID>
<name>OUT</name></connection>
<connection>
<GID>1397</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-502.5,274,-502.5</points>
<connection>
<GID>1391</GID>
<name>OUT</name></connection>
<connection>
<GID>1396</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-506.5,274,-506.5</points>
<connection>
<GID>1392</GID>
<name>OUT</name></connection>
<connection>
<GID>1399</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-510.5,274,-510.5</points>
<connection>
<GID>1393</GID>
<name>OUT</name></connection>
<connection>
<GID>1400</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-514.5,274,-514.5</points>
<connection>
<GID>1394</GID>
<name>OUT</name></connection>
<connection>
<GID>1401</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-518.5,274,-518.5</points>
<connection>
<GID>1395</GID>
<name>OUT</name></connection>
<connection>
<GID>1402</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1110</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>274,-524.5,274,-524.5</points>
<connection>
<GID>1403</GID>
<name>N_in0</name></connection>
<connection>
<GID>1404</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-532.5,274,-532.5</points>
<connection>
<GID>1406</GID>
<name>OUT</name></connection>
<connection>
<GID>1414</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-528.5,274,-528.5</points>
<connection>
<GID>1405</GID>
<name>OUT</name></connection>
<connection>
<GID>1413</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-536.5,274,-536.5</points>
<connection>
<GID>1407</GID>
<name>OUT</name></connection>
<connection>
<GID>1412</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-540.5,274,-540.5</points>
<connection>
<GID>1408</GID>
<name>OUT</name></connection>
<connection>
<GID>1415</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-544.5,274,-544.5</points>
<connection>
<GID>1409</GID>
<name>OUT</name></connection>
<connection>
<GID>1416</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-548.5,274,-548.5</points>
<connection>
<GID>1410</GID>
<name>OUT</name></connection>
<connection>
<GID>1417</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-552.5,274,-552.5</points>
<connection>
<GID>1411</GID>
<name>OUT</name></connection>
<connection>
<GID>1418</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1118</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-517.5,268,-517.5</points>
<connection>
<GID>1395</GID>
<name>IN_0</name></connection>
<connection>
<GID>1425</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-551.5,257,-413</points>
<intersection>-551.5 18</intersection>
<intersection>-547.5 17</intersection>
<intersection>-543.5 16</intersection>
<intersection>-539.5 15</intersection>
<intersection>-535.5 14</intersection>
<intersection>-531.5 13</intersection>
<intersection>-527.5 12</intersection>
<intersection>-523.5 11</intersection>
<intersection>-517.5 2</intersection>
<intersection>-513.5 9</intersection>
<intersection>-509.5 8</intersection>
<intersection>-505.5 7</intersection>
<intersection>-501.5 6</intersection>
<intersection>-497.5 5</intersection>
<intersection>-493.5 4</intersection>
<intersection>-489.5 3</intersection>
<intersection>-482 38</intersection>
<intersection>-478 37</intersection>
<intersection>-474 36</intersection>
<intersection>-470 35</intersection>
<intersection>-466 34</intersection>
<intersection>-462 33</intersection>
<intersection>-458 32</intersection>
<intersection>-454 31</intersection>
<intersection>-448 22</intersection>
<intersection>-444 29</intersection>
<intersection>-440 28</intersection>
<intersection>-436 27</intersection>
<intersection>-432 26</intersection>
<intersection>-428 25</intersection>
<intersection>-424 24</intersection>
<intersection>-420 23</intersection>
<intersection>-413 21</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>257,-517.5,264,-517.5</points>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>257,-489.5,264,-489.5</points>
<connection>
<GID>1388</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>257,-493.5,264,-493.5</points>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>257,-497.5,264,-497.5</points>
<connection>
<GID>1420</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>257,-501.5,264,-501.5</points>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>257,-505.5,264,-505.5</points>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>257,-509.5,264,-509.5</points>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>257,-513.5,264,-513.5</points>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>257,-523.5,268,-523.5</points>
<connection>
<GID>1404</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>257,-527.5,268,-527.5</points>
<connection>
<GID>1405</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>257,-531.5,268,-531.5</points>
<connection>
<GID>1406</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>257,-535.5,268,-535.5</points>
<connection>
<GID>1407</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>257,-539.5,268,-539.5</points>
<connection>
<GID>1408</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>257,-543.5,268,-543.5</points>
<connection>
<GID>1409</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>257,-547.5,268,-547.5</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>257,-551.5,268,-551.5</points>
<connection>
<GID>1411</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>204,-413,257,-413</points>
<intersection>204 40</intersection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>257,-448,264,-448</points>
<connection>
<GID>1384</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>257,-420,264,-420</points>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>257,-424,264,-424</points>
<connection>
<GID>1378</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>257,-428,264,-428</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>257,-432,264,-432</points>
<connection>
<GID>1380</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>257,-436,264,-436</points>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>257,-440,264,-440</points>
<connection>
<GID>1382</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>257,-444,264,-444</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>257,-454,268,-454</points>
<connection>
<GID>1363</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>257,-458,268,-458</points>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>257,-462,268,-462</points>
<connection>
<GID>1365</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>257,-466,268,-466</points>
<connection>
<GID>1366</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>257,-470,268,-470</points>
<connection>
<GID>1367</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>257,-474,268,-474</points>
<connection>
<GID>1368</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>257,-478,268,-478</points>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>257,-482,268,-482</points>
<connection>
<GID>1370</GID>
<name>IN_0</name></connection>
<intersection>257 0</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>204,-466.5,204,-413</points>
<intersection>-466.5 42</intersection>
<intersection>-413 21</intersection></vsegment>
<hsegment>
<ID>42</ID>
<points>202.5,-466.5,204,-466.5</points>
<connection>
<GID>232</GID>
<name>Q</name></connection>
<intersection>204 40</intersection></hsegment></shape></wire>
<wire>
<ID>1120</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-513.5,268,-513.5</points>
<connection>
<GID>1394</GID>
<name>IN_0</name></connection>
<connection>
<GID>1424</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1121</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-509.5,268,-509.5</points>
<connection>
<GID>1393</GID>
<name>IN_0</name></connection>
<connection>
<GID>1423</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1122</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-505.5,268,-505.5</points>
<connection>
<GID>1392</GID>
<name>IN_0</name></connection>
<connection>
<GID>1422</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1123</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-501.5,268,-501.5</points>
<connection>
<GID>1391</GID>
<name>IN_0</name></connection>
<connection>
<GID>1421</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1124</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-497.5,268,-497.5</points>
<connection>
<GID>1390</GID>
<name>IN_0</name></connection>
<connection>
<GID>1420</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1125</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268,-493.5,268,-493.5</points>
<connection>
<GID>1389</GID>
<name>IN_0</name></connection>
<connection>
<GID>1419</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-468,302,-468</points>
<connection>
<GID>1335</GID>
<name>OUT</name></connection>
<connection>
<GID>1434</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-472,302,-472</points>
<connection>
<GID>1336</GID>
<name>OUT</name></connection>
<connection>
<GID>1436</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-496,302,-496</points>
<connection>
<GID>1342</GID>
<name>OUT</name></connection>
<connection>
<GID>1441</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-476,302,-476</points>
<connection>
<GID>1337</GID>
<name>OUT</name></connection>
<connection>
<GID>1437</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-480,302,-480</points>
<connection>
<GID>1338</GID>
<name>OUT</name></connection>
<connection>
<GID>1435</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-484,302,-484</points>
<connection>
<GID>1339</GID>
<name>OUT</name></connection>
<connection>
<GID>1438</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-488,302,-488</points>
<connection>
<GID>1340</GID>
<name>OUT</name></connection>
<connection>
<GID>1439</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-492,302,-492</points>
<connection>
<GID>1341</GID>
<name>OUT</name></connection>
<connection>
<GID>1440</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>1134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300,-431.5,300,-421</points>
<intersection>-431.5 1</intersection>
<intersection>-421 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300,-431.5,302,-431.5</points>
<connection>
<GID>1426</GID>
<name>N_in0</name></connection>
<intersection>300 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-421,300,-421</points>
<connection>
<GID>1345</GID>
<name>N_in1</name></connection>
<intersection>300 0</intersection></hsegment></shape></wire>
<wire>
<ID>1135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-435.5,298.5,-425</points>
<intersection>-435.5 2</intersection>
<intersection>-425 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-425,298.5,-425</points>
<connection>
<GID>1356</GID>
<name>N_in1</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298.5,-435.5,302,-435.5</points>
<connection>
<GID>1428</GID>
<name>N_in0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297,-439.5,297,-429</points>
<intersection>-439.5 2</intersection>
<intersection>-429 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-429,297,-429</points>
<connection>
<GID>1357</GID>
<name>N_in1</name></connection>
<intersection>297 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>297,-439.5,302,-439.5</points>
<connection>
<GID>1429</GID>
<name>N_in0</name></connection>
<intersection>297 0</intersection></hsegment></shape></wire>
<wire>
<ID>1137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,-443.5,295.5,-433</points>
<intersection>-443.5 1</intersection>
<intersection>-433 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,-443.5,302,-443.5</points>
<connection>
<GID>1427</GID>
<name>N_in0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-433,295.5,-433</points>
<connection>
<GID>1355</GID>
<name>N_in1</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294.5,-447.5,294.5,-437</points>
<intersection>-447.5 1</intersection>
<intersection>-437 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294.5,-447.5,302,-447.5</points>
<connection>
<GID>1430</GID>
<name>N_in0</name></connection>
<intersection>294.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-437,294.5,-437</points>
<connection>
<GID>1358</GID>
<name>N_in1</name></connection>
<intersection>294.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-451.5,293,-441</points>
<intersection>-451.5 2</intersection>
<intersection>-441 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-441,293,-441</points>
<connection>
<GID>1359</GID>
<name>N_in1</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>293,-451.5,302,-451.5</points>
<connection>
<GID>1431</GID>
<name>N_in0</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>1140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-455.5,292,-445</points>
<intersection>-455.5 1</intersection>
<intersection>-445 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-455.5,302,-455.5</points>
<connection>
<GID>1432</GID>
<name>N_in0</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-445,292,-445</points>
<connection>
<GID>1360</GID>
<name>N_in1</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>1141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>291,-459.5,291,-449</points>
<intersection>-459.5 2</intersection>
<intersection>-449 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-449,291,-449</points>
<connection>
<GID>1361</GID>
<name>N_in1</name></connection>
<intersection>291 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>291,-459.5,302,-459.5</points>
<connection>
<GID>1433</GID>
<name>N_in0</name></connection>
<intersection>291 0</intersection></hsegment></shape></wire>
<wire>
<ID>1142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289,-467,289,-455</points>
<intersection>-467 1</intersection>
<intersection>-455 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>289,-467,296,-467</points>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection>
<intersection>289 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-455,289,-455</points>
<connection>
<GID>1362</GID>
<name>N_in1</name></connection>
<intersection>289 0</intersection></hsegment></shape></wire>
<wire>
<ID>1143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-471,287.5,-459</points>
<intersection>-471 1</intersection>
<intersection>-459 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287.5,-471,296,-471</points>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection>
<intersection>287.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-459,287.5,-459</points>
<connection>
<GID>1372</GID>
<name>N_in1</name></connection>
<intersection>287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-475,286,-463</points>
<intersection>-475 1</intersection>
<intersection>-463 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-475,296,-475</points>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-463,286,-463</points>
<connection>
<GID>1373</GID>
<name>N_in1</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>1145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-479,284.5,-467</points>
<intersection>-479 1</intersection>
<intersection>-467 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-479,296,-479</points>
<connection>
<GID>1338</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-467,284.5,-467</points>
<connection>
<GID>1371</GID>
<name>N_in1</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283,-483,283,-471</points>
<intersection>-483 1</intersection>
<intersection>-471 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283,-483,296,-483</points>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection>
<intersection>283 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-471,283,-471</points>
<connection>
<GID>1374</GID>
<name>N_in1</name></connection>
<intersection>283 0</intersection></hsegment></shape></wire>
<wire>
<ID>1147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281.5,-487,281.5,-475</points>
<intersection>-487 1</intersection>
<intersection>-475 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-487,296,-487</points>
<connection>
<GID>1340</GID>
<name>IN_0</name></connection>
<intersection>281.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-475,281.5,-475</points>
<connection>
<GID>1375</GID>
<name>N_in1</name></connection>
<intersection>281.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-491,280,-479</points>
<intersection>-491 1</intersection>
<intersection>-479 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280,-491,296,-491</points>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-479,280,-479</points>
<connection>
<GID>1376</GID>
<name>N_in1</name></connection>
<intersection>280 0</intersection></hsegment></shape></wire>
<wire>
<ID>1149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-495,278.5,-483</points>
<intersection>-495 1</intersection>
<intersection>-483 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278.5,-495,296,-495</points>
<connection>
<GID>1342</GID>
<name>IN_0</name></connection>
<intersection>278.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-483,278.5,-483</points>
<connection>
<GID>1377</GID>
<name>N_in1</name></connection>
<intersection>278.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-490.5,290,-469</points>
<intersection>-490.5 2</intersection>
<intersection>-469 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-469,296,-469</points>
<connection>
<GID>1335</GID>
<name>IN_1</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-490.5,290,-490.5</points>
<connection>
<GID>1386</GID>
<name>N_in1</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>1151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-494.5,288.5,-473</points>
<intersection>-494.5 1</intersection>
<intersection>-473 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-494.5,288.5,-494.5</points>
<connection>
<GID>1397</GID>
<name>N_in1</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288.5,-473,296,-473</points>
<connection>
<GID>1336</GID>
<name>IN_1</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-498.5,287,-477</points>
<intersection>-498.5 1</intersection>
<intersection>-477 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-498.5,287,-498.5</points>
<connection>
<GID>1398</GID>
<name>N_in1</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287,-477,296,-477</points>
<connection>
<GID>1337</GID>
<name>IN_1</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire>
<wire>
<ID>1153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-502.5,285.5,-481</points>
<intersection>-502.5 1</intersection>
<intersection>-481 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-502.5,285.5,-502.5</points>
<connection>
<GID>1396</GID>
<name>N_in1</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-481,296,-481</points>
<connection>
<GID>1338</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-506.5,284,-485</points>
<intersection>-506.5 1</intersection>
<intersection>-485 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-506.5,284,-506.5</points>
<connection>
<GID>1399</GID>
<name>N_in1</name></connection>
<intersection>284 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>284,-485,296,-485</points>
<connection>
<GID>1339</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment></shape></wire>
<wire>
<ID>1155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282.5,-510.5,282.5,-489</points>
<intersection>-510.5 1</intersection>
<intersection>-489 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-510.5,282.5,-510.5</points>
<connection>
<GID>1400</GID>
<name>N_in1</name></connection>
<intersection>282.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>282.5,-489,296,-489</points>
<connection>
<GID>1340</GID>
<name>IN_1</name></connection>
<intersection>282.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-514.5,281,-493</points>
<intersection>-514.5 1</intersection>
<intersection>-493 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-514.5,281,-514.5</points>
<connection>
<GID>1401</GID>
<name>N_in1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281,-493,296,-493</points>
<connection>
<GID>1341</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>1157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-518.5,279.5,-497</points>
<intersection>-518.5 1</intersection>
<intersection>-497 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-518.5,279.5,-518.5</points>
<connection>
<GID>1402</GID>
<name>N_in1</name></connection>
<intersection>279.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>279.5,-497,296,-497</points>
<connection>
<GID>1342</GID>
<name>IN_1</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-524.5,286.5,-508</points>
<intersection>-524.5 2</intersection>
<intersection>-508 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286.5,-508,302.5,-508</points>
<connection>
<GID>1324</GID>
<name>N_in0</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-524.5,286.5,-524.5</points>
<connection>
<GID>1403</GID>
<name>N_in1</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-528.5,288.5,-512</points>
<intersection>-528.5 2</intersection>
<intersection>-512 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-512,302.5,-512</points>
<connection>
<GID>1326</GID>
<name>N_in0</name></connection>
<intersection>288.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-528.5,288.5,-528.5</points>
<connection>
<GID>1413</GID>
<name>N_in1</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-532.5,290,-516</points>
<intersection>-532.5 2</intersection>
<intersection>-516 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>290,-516,302.5,-516</points>
<connection>
<GID>1327</GID>
<name>N_in0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-532.5,290,-532.5</points>
<connection>
<GID>1414</GID>
<name>N_in1</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>1161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>292,-536.5,292,-520</points>
<intersection>-536.5 2</intersection>
<intersection>-520 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292,-520,302.5,-520</points>
<connection>
<GID>1325</GID>
<name>N_in0</name></connection>
<intersection>292 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-536.5,292,-536.5</points>
<connection>
<GID>1412</GID>
<name>N_in1</name></connection>
<intersection>292 0</intersection></hsegment></shape></wire>
<wire>
<ID>1162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-540.5,294,-524</points>
<intersection>-540.5 2</intersection>
<intersection>-524 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>294,-524,302.5,-524</points>
<connection>
<GID>1328</GID>
<name>N_in0</name></connection>
<intersection>294 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-540.5,294,-540.5</points>
<connection>
<GID>1415</GID>
<name>N_in1</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>1163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>296.5,-544.5,296.5,-528</points>
<intersection>-544.5 2</intersection>
<intersection>-528 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>296.5,-528,302.5,-528</points>
<connection>
<GID>1329</GID>
<name>N_in0</name></connection>
<intersection>296.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-544.5,296.5,-544.5</points>
<connection>
<GID>1416</GID>
<name>N_in1</name></connection>
<intersection>296.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-548.5,298.5,-532</points>
<intersection>-548.5 1</intersection>
<intersection>-532 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-548.5,298.5,-548.5</points>
<connection>
<GID>1417</GID>
<name>N_in1</name></connection>
<intersection>298.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>298.5,-532,302.5,-532</points>
<connection>
<GID>1330</GID>
<name>N_in0</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>300.5,-552.5,300.5,-536</points>
<intersection>-552.5 2</intersection>
<intersection>-536 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>300.5,-536,302.5,-536</points>
<connection>
<GID>1331</GID>
<name>N_in0</name></connection>
<intersection>300.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>276,-552.5,300.5,-552.5</points>
<connection>
<GID>1418</GID>
<name>N_in1</name></connection>
<intersection>300.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-423,243,-423</points>
<connection>
<GID>1464</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1479</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-427,243,-427</points>
<connection>
<GID>1466</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1480</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-431,243,-431</points>
<connection>
<GID>1468</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1481</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-435,243,-435</points>
<connection>
<GID>1470</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1482</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-439,243,-439</points>
<connection>
<GID>1472</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1483</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-443,243,-443</points>
<connection>
<GID>1474</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1484</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-447,243,-447</points>
<connection>
<GID>1476</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1485</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>243,-451,243,-451</points>
<connection>
<GID>1478</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1486</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>231,-421,243,-421</points>
<connection>
<GID>1479</GID>
<name>IN_0</name></connection>
<connection>
<GID>1487</GID>
<name>OUT_0</name></connection>
<intersection>231 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>231,-449,231,-421</points>
<intersection>-449 4</intersection>
<intersection>-445 10</intersection>
<intersection>-441 9</intersection>
<intersection>-437 8</intersection>
<intersection>-433 7</intersection>
<intersection>-429 6</intersection>
<intersection>-425 5</intersection>
<intersection>-421 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>231,-449,243,-449</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>231,-425,243,-425</points>
<connection>
<GID>1480</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>231,-429,243,-429</points>
<connection>
<GID>1481</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>231,-433,243,-433</points>
<connection>
<GID>1482</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>231,-437,243,-437</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>231,-441,243,-441</points>
<connection>
<GID>1484</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>231,-445,243,-445</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<intersection>231 3</intersection></hsegment></shape></wire>
<wire>
<ID>1193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>179.5,-462.5,236.5,-462.5</points>
<intersection>179.5 12</intersection>
<intersection>236.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236.5,-518.5,236.5,-462.5</points>
<intersection>-518.5 4</intersection>
<intersection>-514.5 10</intersection>
<intersection>-510.5 9</intersection>
<intersection>-506.5 8</intersection>
<intersection>-502.5 7</intersection>
<intersection>-498.5 6</intersection>
<intersection>-494.5 5</intersection>
<intersection>-490.5 28</intersection>
<intersection>-462.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>236.5,-518.5,242.5,-518.5</points>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>236.5,-494.5,242.5,-494.5</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>236.5,-498.5,242.5,-498.5</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>236.5,-502.5,242.5,-502.5</points>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>236.5,-506.5,242.5,-506.5</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>236.5,-510.5,242.5,-510.5</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>236.5,-514.5,242.5,-514.5</points>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>179.5,-466.5,179.5,-421</points>
<connection>
<GID>231</GID>
<name>Q</name></connection>
<intersection>-463.5 21</intersection>
<intersection>-462.5 1</intersection>
<intersection>-421 26</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>179.5,-463.5,180.5,-463.5</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>179.5 12</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>179.5,-421,227,-421</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<intersection>179.5 12</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>236.5,-490.5,242.5,-490.5</points>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection>
<intersection>236.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,-533,325,-526</points>
<connection>
<GID>1507</GID>
<name>clock</name></connection>
<intersection>-533 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-533,325,-533</points>
<connection>
<GID>1508</GID>
<name>CLK</name></connection>
<intersection>325 0</intersection></hsegment></shape></wire>
<wire>
<ID>1203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-455.5,321,-452.5</points>
<connection>
<GID>1506</GID>
<name>clock</name></connection>
<intersection>-455.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>320,-455.5,321,-455.5</points>
<connection>
<GID>1509</GID>
<name>CLK</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>1204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-441.5,321,-440.5</points>
<connection>
<GID>1506</GID>
<name>load</name></connection>
<intersection>-440.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-440.5,321,-440.5</points>
<connection>
<GID>1510</GID>
<name>OUT_0</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>1205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-489.5,323,-484.5</points>
<connection>
<GID>1511</GID>
<name>clock</name></connection>
<intersection>-489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321,-489.5,323,-489.5</points>
<connection>
<GID>1512</GID>
<name>CLK</name></connection>
<intersection>323 0</intersection></hsegment></shape></wire>
<wire>
<ID>1206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-473.5,323,-472</points>
<connection>
<GID>1511</GID>
<name>load</name></connection>
<intersection>-472 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322.5,-472,323,-472</points>
<connection>
<GID>1513</GID>
<name>OUT_0</name></connection>
<intersection>323 0</intersection></hsegment></shape></wire>
<wire>
<ID>1207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,-515,325,-511</points>
<connection>
<GID>1507</GID>
<name>load</name></connection>
<intersection>-511 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323.5,-511,325,-511</points>
<connection>
<GID>1514</GID>
<name>OUT_0</name></connection>
<intersection>325 0</intersection></hsegment></shape></wire>
<wire>
<ID>1208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101.5,74,110,74</points>
<connection>
<GID>1515</GID>
<name>J</name></connection>
<intersection>101.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>101.5,65,101.5,74</points>
<connection>
<GID>1521</GID>
<name>carry_out</name></connection>
<intersection>70 5</intersection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>101.5,70,110,70</points>
<connection>
<GID>1515</GID>
<name>K</name></connection>
<intersection>101.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,65,99.5,65</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1521</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>1212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,65,100.5,71</points>
<connection>
<GID>1521</GID>
<name>count_up</name></connection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,71,100.5,71</points>
<intersection>75 2</intersection>
<intersection>100.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,54.5,75,71</points>
<intersection>54.5 3</intersection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>69,54.5,75,54.5</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-18.5,295.5,-18.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<connection>
<GID>656</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>285,-54.5,285,-20.5</points>
<intersection>-54.5 19</intersection>
<intersection>-27 23</intersection>
<intersection>-20.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>285,-20.5,295.5,-20.5</points>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<intersection>285 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>285,-54.5,295.5,-54.5</points>
<connection>
<GID>672</GID>
<name>IN_1</name></connection>
<intersection>285 3</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>282,-27,285,-27</points>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection>
<intersection>285 3</intersection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-19.5,301.5,-19.5</points>
<connection>
<GID>654</GID>
<name>N_in0</name></connection>
<connection>
<GID>655</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-58.5,285.5,-24.5</points>
<intersection>-58.5 3</intersection>
<intersection>-29 6</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285.5,-24.5,295.5,-24.5</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>285.5,-58.5,295.5,-58.5</points>
<connection>
<GID>673</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>282,-29,285.5,-29</points>
<connection>
<GID>646</GID>
<name>OUT_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-62.5,286,-28.5</points>
<intersection>-62.5 3</intersection>
<intersection>-31 6</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-28.5,295.5,-28.5</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286,-62.5,295.5,-62.5</points>
<connection>
<GID>674</GID>
<name>IN_1</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>282,-31,286,-31</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>286.5,-66.5,286.5,-32.5</points>
<intersection>-66.5 5</intersection>
<intersection>-33 11</intersection>
<intersection>-32.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>286.5,-66.5,295.5,-66.5</points>
<connection>
<GID>675</GID>
<name>IN_1</name></connection>
<intersection>286.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>286.5,-32.5,295.5,-32.5</points>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<intersection>286.5 4</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>282,-33,286.5,-33</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<intersection>286.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>287,-70.5,287,-35</points>
<intersection>-70.5 4</intersection>
<intersection>-36.5 8</intersection>
<intersection>-35 11</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287,-70.5,295.5,-70.5</points>
<connection>
<GID>676</GID>
<name>IN_1</name></connection>
<intersection>287 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>287,-36.5,295.5,-36.5</points>
<connection>
<GID>660</GID>
<name>IN_1</name></connection>
<intersection>287 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>282,-35,287,-35</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<intersection>287 3</intersection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>282,-37,295.5,-37</points>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<intersection>287.5 3</intersection>
<intersection>295.5 11</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>287.5,-74.5,287.5,-37</points>
<intersection>-74.5 4</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,-74.5,295.5,-74.5</points>
<connection>
<GID>677</GID>
<name>IN_1</name></connection>
<intersection>287.5 3</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>295.5,-40.5,295.5,-37</points>
<connection>
<GID>661</GID>
<name>IN_1</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>288,-44.5,295.5,-44.5</points>
<connection>
<GID>662</GID>
<name>IN_1</name></connection>
<intersection>288 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,-78.5,288,-39</points>
<intersection>-78.5 4</intersection>
<intersection>-44.5 1</intersection>
<intersection>-39 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,-78.5,295.5,-78.5</points>
<connection>
<GID>678</GID>
<name>IN_1</name></connection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>282,-39,288,-39</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>288.5,-82.5,288.5,-41</points>
<intersection>-82.5 4</intersection>
<intersection>-48.5 5</intersection>
<intersection>-41 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,-82.5,295.5,-82.5</points>
<connection>
<GID>679</GID>
<name>IN_1</name></connection>
<intersection>288.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>288.5,-48.5,295.5,-48.5</points>
<connection>
<GID>663</GID>
<name>IN_1</name></connection>
<intersection>288.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>282,-41,288.5,-41</points>
<connection>
<GID>652</GID>
<name>OUT_0</name></connection>
<intersection>288.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-27.5,301.5,-27.5</points>
<connection>
<GID>658</GID>
<name>OUT</name></connection>
<connection>
<GID>666</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-23.5,301.5,-23.5</points>
<connection>
<GID>657</GID>
<name>OUT</name></connection>
<connection>
<GID>665</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-31.5,301.5,-31.5</points>
<connection>
<GID>659</GID>
<name>OUT</name></connection>
<connection>
<GID>664</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-35.5,301.5,-35.5</points>
<connection>
<GID>660</GID>
<name>OUT</name></connection>
<connection>
<GID>667</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-39.5,301.5,-39.5</points>
<connection>
<GID>661</GID>
<name>OUT</name></connection>
<connection>
<GID>668</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-43.5,301.5,-43.5</points>
<connection>
<GID>662</GID>
<name>OUT</name></connection>
<connection>
<GID>669</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-47.5,301.5,-47.5</points>
<connection>
<GID>663</GID>
<name>OUT</name></connection>
<connection>
<GID>670</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-53.5,301.5,-53.5</points>
<connection>
<GID>671</GID>
<name>N_in0</name></connection>
<connection>
<GID>672</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-61.5,301.5,-61.5</points>
<connection>
<GID>674</GID>
<name>OUT</name></connection>
<connection>
<GID>682</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-57.5,301.5,-57.5</points>
<connection>
<GID>673</GID>
<name>OUT</name></connection>
<connection>
<GID>681</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-65.5,301.5,-65.5</points>
<connection>
<GID>675</GID>
<name>OUT</name></connection>
<connection>
<GID>680</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-69.5,301.5,-69.5</points>
<connection>
<GID>676</GID>
<name>OUT</name></connection>
<connection>
<GID>683</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-73.5,301.5,-73.5</points>
<connection>
<GID>677</GID>
<name>OUT</name></connection>
<connection>
<GID>684</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-77.5,301.5,-77.5</points>
<connection>
<GID>678</GID>
<name>OUT</name></connection>
<connection>
<GID>685</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-81.5,301.5,-81.5</points>
<connection>
<GID>679</GID>
<name>OUT</name></connection>
<connection>
<GID>686</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-46.5,295.5,-46.5</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-42.5,295.5,-42.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<connection>
<GID>692</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-38.5,295.5,-38.5</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-34.5,295.5,-34.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-30.5,295.5,-30.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<connection>
<GID>689</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-26.5,295.5,-26.5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<connection>
<GID>688</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-22.5,295.5,-22.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-88,295.5,-88</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<connection>
<GID>699</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-96.5,285,-96.5</points>
<connection>
<GID>696</GID>
<name>OUT_0</name></connection>
<intersection>285 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>285,-124,285,-90</points>
<intersection>-124 19</intersection>
<intersection>-96.5 1</intersection>
<intersection>-90 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>285,-90,295.5,-90</points>
<connection>
<GID>698</GID>
<name>IN_1</name></connection>
<intersection>285 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>285,-124,295.5,-124</points>
<connection>
<GID>722</GID>
<name>IN_1</name></connection>
<intersection>285 3</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-89,301.5,-89</points>
<connection>
<GID>697</GID>
<name>N_in0</name></connection>
<connection>
<GID>698</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-128,285.5,-94</points>
<intersection>-128 3</intersection>
<intersection>-98.5 2</intersection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>285.5,-94,295.5,-94</points>
<connection>
<GID>707</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-98.5,285.5,-98.5</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>285.5,-128,295.5,-128</points>
<connection>
<GID>723</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-132,286,-98</points>
<intersection>-132 3</intersection>
<intersection>-100.5 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-98,295.5,-98</points>
<connection>
<GID>708</GID>
<name>IN_1</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-100.5,286,-100.5</points>
<connection>
<GID>701</GID>
<name>OUT_0</name></connection>
<intersection>286 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286,-132,295.5,-132</points>
<connection>
<GID>724</GID>
<name>IN_1</name></connection>
<intersection>286 0</intersection></hsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-102.5,286.5,-102.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>286.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>286.5,-136,286.5,-102</points>
<intersection>-136 5</intersection>
<intersection>-102.5 1</intersection>
<intersection>-102 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>286.5,-136,295.5,-136</points>
<connection>
<GID>725</GID>
<name>IN_1</name></connection>
<intersection>286.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>286.5,-102,295.5,-102</points>
<connection>
<GID>709</GID>
<name>IN_1</name></connection>
<intersection>286.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-104.5,287,-104.5</points>
<connection>
<GID>703</GID>
<name>OUT_0</name></connection>
<intersection>287 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>287,-140,287,-104.5</points>
<intersection>-140 4</intersection>
<intersection>-106 8</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287,-140,295.5,-140</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<intersection>287 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>287,-106,295.5,-106</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<intersection>287 3</intersection></hsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-106.5,287.5,-106.5</points>
<connection>
<GID>704</GID>
<name>OUT_0</name></connection>
<intersection>287.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>287.5,-144,287.5,-106.5</points>
<intersection>-144 4</intersection>
<intersection>-110 8</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>287.5,-144,295.5,-144</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<intersection>287.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>287.5,-110,295.5,-110</points>
<connection>
<GID>711</GID>
<name>IN_1</name></connection>
<intersection>287.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286,-114,286,-108.5</points>
<intersection>-114 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>286,-114,295.5,-114</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>286 0</intersection>
<intersection>288 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>281.5,-108.5,286,-108.5</points>
<connection>
<GID>705</GID>
<name>OUT_0</name></connection>
<intersection>286 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288,-148,288,-114</points>
<intersection>-148 4</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288,-148,295.5,-148</points>
<connection>
<GID>728</GID>
<name>IN_1</name></connection>
<intersection>288 3</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-110.5,288.5,-110.5</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>288.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>288.5,-152,288.5,-110.5</points>
<intersection>-152 4</intersection>
<intersection>-118 5</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>288.5,-152,295.5,-152</points>
<connection>
<GID>729</GID>
<name>IN_1</name></connection>
<intersection>288.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>288.5,-118,295.5,-118</points>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>288.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-97,301.5,-97</points>
<connection>
<GID>708</GID>
<name>OUT</name></connection>
<connection>
<GID>716</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-93,301.5,-93</points>
<connection>
<GID>707</GID>
<name>OUT</name></connection>
<connection>
<GID>715</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-101,301.5,-101</points>
<connection>
<GID>709</GID>
<name>OUT</name></connection>
<connection>
<GID>714</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-105,301.5,-105</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<connection>
<GID>717</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-109,301.5,-109</points>
<connection>
<GID>711</GID>
<name>OUT</name></connection>
<connection>
<GID>718</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-113,301.5,-113</points>
<connection>
<GID>712</GID>
<name>OUT</name></connection>
<connection>
<GID>719</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-117,301.5,-117</points>
<connection>
<GID>713</GID>
<name>OUT</name></connection>
<connection>
<GID>720</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>301.5,-123,301.5,-123</points>
<connection>
<GID>721</GID>
<name>N_in0</name></connection>
<connection>
<GID>722</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-131,301.5,-131</points>
<connection>
<GID>724</GID>
<name>OUT</name></connection>
<connection>
<GID>732</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-127,301.5,-127</points>
<connection>
<GID>723</GID>
<name>OUT</name></connection>
<connection>
<GID>731</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-135,301.5,-135</points>
<connection>
<GID>725</GID>
<name>OUT</name></connection>
<connection>
<GID>730</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-139,301.5,-139</points>
<connection>
<GID>726</GID>
<name>OUT</name></connection>
<connection>
<GID>733</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-143,301.5,-143</points>
<connection>
<GID>727</GID>
<name>OUT</name></connection>
<connection>
<GID>734</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-147,301.5,-147</points>
<connection>
<GID>728</GID>
<name>OUT</name></connection>
<connection>
<GID>735</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-151,301.5,-151</points>
<connection>
<GID>729</GID>
<name>OUT</name></connection>
<connection>
<GID>736</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-116,295.5,-116</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<connection>
<GID>743</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284.5,-150,284.5,-11.5</points>
<intersection>-150 18</intersection>
<intersection>-146 17</intersection>
<intersection>-142 16</intersection>
<intersection>-138 15</intersection>
<intersection>-134 14</intersection>
<intersection>-130 13</intersection>
<intersection>-126 12</intersection>
<intersection>-122 11</intersection>
<intersection>-116 2</intersection>
<intersection>-112 9</intersection>
<intersection>-108 8</intersection>
<intersection>-104 7</intersection>
<intersection>-100 6</intersection>
<intersection>-96 5</intersection>
<intersection>-92 4</intersection>
<intersection>-88 3</intersection>
<intersection>-80.5 38</intersection>
<intersection>-76.5 37</intersection>
<intersection>-72.5 36</intersection>
<intersection>-68.5 35</intersection>
<intersection>-64.5 34</intersection>
<intersection>-60.5 33</intersection>
<intersection>-56.5 32</intersection>
<intersection>-52.5 31</intersection>
<intersection>-46.5 22</intersection>
<intersection>-42.5 29</intersection>
<intersection>-38.5 28</intersection>
<intersection>-34.5 27</intersection>
<intersection>-30.5 26</intersection>
<intersection>-26.5 25</intersection>
<intersection>-22.5 24</intersection>
<intersection>-18.5 23</intersection>
<intersection>-11.5 21</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>284.5,-116,291.5,-116</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>284.5,-88,291.5,-88</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>284.5,-92,291.5,-92</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>284.5,-96,291.5,-96</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>284.5,-100,291.5,-100</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>284.5,-104,291.5,-104</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>284.5,-108,291.5,-108</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>284.5,-112,291.5,-112</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>284.5,-122,295.5,-122</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>284.5,-126,295.5,-126</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>284.5,-130,295.5,-130</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>284.5,-134,295.5,-134</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>284.5,-138,295.5,-138</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>284.5,-142,295.5,-142</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>284.5,-146,295.5,-146</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>284.5,-150,295.5,-150</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>272,-11.5,284.5,-11.5</points>
<connection>
<GID>653</GID>
<name>OUT_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>284.5,-46.5,291.5,-46.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>284.5,-18.5,291.5,-18.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>284.5,-22.5,291.5,-22.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>284.5,-26.5,291.5,-26.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>284.5,-30.5,291.5,-30.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>284.5,-34.5,291.5,-34.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>284.5,-38.5,291.5,-38.5</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>284.5,-42.5,291.5,-42.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>284.5,-52.5,295.5,-52.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>284.5,-56.5,295.5,-56.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>284.5,-60.5,295.5,-60.5</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>284.5,-64.5,295.5,-64.5</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>284.5,-68.5,295.5,-68.5</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>284.5,-72.5,295.5,-72.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>284.5,-76.5,295.5,-76.5</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>284.5,-80.5,295.5,-80.5</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>284.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-112,295.5,-112</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<connection>
<GID>742</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-108,295.5,-108</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<connection>
<GID>741</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-104,295.5,-104</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-100,295.5,-100</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-96,295.5,-96</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-92,295.5,-92</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-29,278,-29</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-27,278,-27</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<connection>
<GID>745</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-35,278,-35</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-37,278,-37</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<connection>
<GID>750</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-31,278,-31</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-41,278,-41</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-39,278,-39</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-33,278,-33</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-66.5,329.5,-66.5</points>
<connection>
<GID>780</GID>
<name>OUT</name></connection>
<connection>
<GID>761</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-70.5,329.5,-70.5</points>
<connection>
<GID>781</GID>
<name>OUT</name></connection>
<connection>
<GID>763</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-94.5,329.5,-94.5</points>
<connection>
<GID>787</GID>
<name>OUT</name></connection>
<connection>
<GID>768</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-74.5,329.5,-74.5</points>
<connection>
<GID>782</GID>
<name>OUT</name></connection>
<connection>
<GID>764</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-78.5,329.5,-78.5</points>
<connection>
<GID>783</GID>
<name>OUT</name></connection>
<connection>
<GID>762</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-82.5,329.5,-82.5</points>
<connection>
<GID>784</GID>
<name>OUT</name></connection>
<connection>
<GID>765</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-86.5,329.5,-86.5</points>
<connection>
<GID>785</GID>
<name>OUT</name></connection>
<connection>
<GID>766</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>329.5,-90.5,329.5,-90.5</points>
<connection>
<GID>786</GID>
<name>OUT</name></connection>
<connection>
<GID>767</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327.5,-30,327.5,-19.5</points>
<intersection>-30 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>327.5,-30,329.5,-30</points>
<connection>
<GID>753</GID>
<name>N_in0</name></connection>
<intersection>327.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-19.5,327.5,-19.5</points>
<connection>
<GID>654</GID>
<name>N_in1</name></connection>
<intersection>327.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,-34,326,-23.5</points>
<intersection>-34 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-23.5,326,-23.5</points>
<connection>
<GID>665</GID>
<name>N_in1</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>326,-34,329.5,-34</points>
<connection>
<GID>755</GID>
<name>N_in0</name></connection>
<intersection>326 0</intersection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-38,324.5,-27.5</points>
<intersection>-38 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-27.5,324.5,-27.5</points>
<connection>
<GID>666</GID>
<name>N_in1</name></connection>
<intersection>324.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>324.5,-38,329.5,-38</points>
<connection>
<GID>756</GID>
<name>N_in0</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>323,-42,323,-31.5</points>
<intersection>-42 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>323,-42,329.5,-42</points>
<connection>
<GID>754</GID>
<name>N_in0</name></connection>
<intersection>323 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-31.5,323,-31.5</points>
<connection>
<GID>664</GID>
<name>N_in1</name></connection>
<intersection>323 0</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322,-46,322,-35.5</points>
<intersection>-46 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>322,-46,329.5,-46</points>
<connection>
<GID>757</GID>
<name>N_in0</name></connection>
<intersection>322 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-35.5,322,-35.5</points>
<connection>
<GID>667</GID>
<name>N_in1</name></connection>
<intersection>322 0</intersection></hsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-50,320.5,-39.5</points>
<intersection>-50 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-39.5,320.5,-39.5</points>
<connection>
<GID>668</GID>
<name>N_in1</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320.5,-50,329.5,-50</points>
<connection>
<GID>758</GID>
<name>N_in0</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-54,319.5,-43.5</points>
<intersection>-54 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-54,329.5,-54</points>
<connection>
<GID>759</GID>
<name>N_in0</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-43.5,319.5,-43.5</points>
<connection>
<GID>669</GID>
<name>N_in1</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-58,318.5,-47.5</points>
<intersection>-58 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-47.5,318.5,-47.5</points>
<connection>
<GID>670</GID>
<name>N_in1</name></connection>
<intersection>318.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>318.5,-58,329.5,-58</points>
<connection>
<GID>760</GID>
<name>N_in0</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317,-65.5,317,-53.5</points>
<intersection>-65.5 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317,-65.5,323.5,-65.5</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>317 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-53.5,317,-53.5</points>
<connection>
<GID>671</GID>
<name>N_in1</name></connection>
<intersection>317 0</intersection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,-69.5,315.5,-57.5</points>
<intersection>-69.5 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315.5,-69.5,323.5,-69.5</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>315.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-57.5,315.5,-57.5</points>
<connection>
<GID>681</GID>
<name>N_in1</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-73.5,314,-61.5</points>
<intersection>-73.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-73.5,323.5,-73.5</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-61.5,314,-61.5</points>
<connection>
<GID>682</GID>
<name>N_in1</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-77.5,313.5,-65.5</points>
<intersection>-77.5 1</intersection>
<intersection>-65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>313.5,-77.5,323.5,-77.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-65.5,313.5,-65.5</points>
<connection>
<GID>680</GID>
<name>N_in1</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-81.5,312.5,-69.5</points>
<intersection>-81.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>312.5,-81.5,323.5,-81.5</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-69.5,312.5,-69.5</points>
<connection>
<GID>683</GID>
<name>N_in1</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-85.5,311,-73.5</points>
<intersection>-85.5 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-85.5,323.5,-85.5</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>311 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-73.5,311,-73.5</points>
<connection>
<GID>684</GID>
<name>N_in1</name></connection>
<intersection>311 0</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>310,-89.5,310,-77.5</points>
<intersection>-89.5 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>310,-89.5,323.5,-89.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>310 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-77.5,310,-77.5</points>
<connection>
<GID>685</GID>
<name>N_in1</name></connection>
<intersection>310 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-93.5,309,-81.5</points>
<intersection>-93.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-93.5,323.5,-93.5</points>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>309 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-81.5,309,-81.5</points>
<connection>
<GID>686</GID>
<name>N_in1</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-89,317.5,-67.5</points>
<intersection>-89 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-67.5,323.5,-67.5</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>317.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-89,317.5,-89</points>
<connection>
<GID>697</GID>
<name>N_in1</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,-93,315.5,-71.5</points>
<intersection>-93 1</intersection>
<intersection>-71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-93,315.5,-93</points>
<connection>
<GID>715</GID>
<name>N_in1</name></connection>
<intersection>315.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>315.5,-71.5,323.5,-71.5</points>
<connection>
<GID>781</GID>
<name>IN_1</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-97,314,-75.5</points>
<intersection>-97 1</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-97,314,-97</points>
<connection>
<GID>716</GID>
<name>N_in1</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>314,-75.5,323.5,-75.5</points>
<connection>
<GID>782</GID>
<name>IN_1</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>313.5,-101,313.5,-79.5</points>
<intersection>-101 1</intersection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-101,313.5,-101</points>
<connection>
<GID>714</GID>
<name>N_in1</name></connection>
<intersection>313.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>313.5,-79.5,323.5,-79.5</points>
<connection>
<GID>783</GID>
<name>IN_1</name></connection>
<intersection>313.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>312.5,-105,312.5,-83.5</points>
<intersection>-105 1</intersection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-105,312.5,-105</points>
<connection>
<GID>717</GID>
<name>N_in1</name></connection>
<intersection>312.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>312.5,-83.5,323.5,-83.5</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>312.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>308,-109,308,-87.5</points>
<intersection>-109 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-109,308,-109</points>
<connection>
<GID>718</GID>
<name>N_in1</name></connection>
<intersection>308 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>308,-87.5,323.5,-87.5</points>
<connection>
<GID>785</GID>
<name>IN_1</name></connection>
<intersection>308 0</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306.5,-113,306.5,-91.5</points>
<intersection>-113 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-113,306.5,-113</points>
<connection>
<GID>719</GID>
<name>N_in1</name></connection>
<intersection>306.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>306.5,-91.5,323.5,-91.5</points>
<connection>
<GID>786</GID>
<name>IN_1</name></connection>
<intersection>306.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>305.5,-117,305.5,-95.5</points>
<intersection>-117 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-117,305.5,-117</points>
<connection>
<GID>720</GID>
<name>N_in1</name></connection>
<intersection>305.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>305.5,-95.5,323.5,-95.5</points>
<connection>
<GID>787</GID>
<name>IN_1</name></connection>
<intersection>305.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>314,-123,314,-106.5</points>
<intersection>-123 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>314,-106.5,330,-106.5</points>
<connection>
<GID>769</GID>
<name>N_in0</name></connection>
<intersection>314 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-123,314,-123</points>
<connection>
<GID>721</GID>
<name>N_in1</name></connection>
<intersection>314 0</intersection></hsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316,-127,316,-110.5</points>
<intersection>-127 2</intersection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>316,-110.5,330,-110.5</points>
<connection>
<GID>771</GID>
<name>N_in0</name></connection>
<intersection>316 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-127,316,-127</points>
<connection>
<GID>731</GID>
<name>N_in1</name></connection>
<intersection>316 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-131,317.5,-114.5</points>
<intersection>-131 2</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-114.5,330,-114.5</points>
<connection>
<GID>772</GID>
<name>N_in0</name></connection>
<intersection>317.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-131,317.5,-131</points>
<connection>
<GID>732</GID>
<name>N_in1</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-135,319.5,-118.5</points>
<intersection>-135 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-118.5,330,-118.5</points>
<connection>
<GID>770</GID>
<name>N_in0</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-135,319.5,-135</points>
<connection>
<GID>730</GID>
<name>N_in1</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321.5,-139,321.5,-122.5</points>
<intersection>-139 2</intersection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>321.5,-122.5,330,-122.5</points>
<connection>
<GID>773</GID>
<name>N_in0</name></connection>
<intersection>321.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-139,321.5,-139</points>
<connection>
<GID>733</GID>
<name>N_in1</name></connection>
<intersection>321.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324,-143,324,-126.5</points>
<intersection>-143 2</intersection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324,-126.5,330,-126.5</points>
<connection>
<GID>774</GID>
<name>N_in0</name></connection>
<intersection>324 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-143,324,-143</points>
<connection>
<GID>734</GID>
<name>N_in1</name></connection>
<intersection>324 0</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>326,-147,326,-130.5</points>
<intersection>-147 1</intersection>
<intersection>-130.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,-147,326,-147</points>
<connection>
<GID>735</GID>
<name>N_in1</name></connection>
<intersection>326 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>326,-130.5,330,-130.5</points>
<connection>
<GID>775</GID>
<name>N_in0</name></connection>
<intersection>326 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>328,-151,328,-134.5</points>
<intersection>-151 2</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>328,-134.5,330,-134.5</points>
<connection>
<GID>776</GID>
<name>N_in0</name></connection>
<intersection>328 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303.5,-151,328,-151</points>
<connection>
<GID>736</GID>
<name>N_in1</name></connection>
<intersection>328 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>146.421,1283.2,1540.42,581.202</PageViewport></page 2>
<page 3>
<PageViewport>-118.962,1678.39,1275.04,976.39</PageViewport></page 3>
<page 4>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 4>
<page 5>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 5>
<page 6>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 6>
<page 7>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 7>
<page 8>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 8>
<page 9>
<PageViewport>0,2797.59,1394,2095.59</PageViewport></page 9></circuit>