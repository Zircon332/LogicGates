<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-225.591,170.048,157.039,-27.2926</PageViewport>
<gate>
<ID>769</ID>
<type>AE_OR2</type>
<position>4,-457.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>770</ID>
<type>AE_OR2</type>
<position>4,-461.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>605 </input>
<output>
<ID>OUT</ID>678 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1</ID>
<type>AE_FULLADDER_4BIT</type>
<position>29.5,-37</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_B_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>96 </output>
<output>
<ID>OUT_3</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_SMALL_INVERTER</type>
<position>3.5,-27</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>772</ID>
<type>AE_REGISTER8</type>
<position>40,-481</position>
<input>
<ID>IN_0</ID>767 </input>
<input>
<ID>IN_1</ID>766 </input>
<input>
<ID>IN_2</ID>765 </input>
<input>
<ID>IN_3</ID>764 </input>
<input>
<ID>IN_4</ID>763 </input>
<input>
<ID>IN_5</ID>762 </input>
<input>
<ID>IN_6</ID>761 </input>
<input>
<ID>IN_7</ID>760 </input>
<input>
<ID>clock</ID>758 </input>
<input>
<ID>load</ID>759 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-27</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>773</ID>
<type>BB_CLOCK</type>
<position>39,-490</position>
<output>
<ID>CLK</ID>758 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,-27</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>27.5,-27</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>34.5,-31</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>-32,23.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>-76,-34</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>-76,-36</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>-76,-38</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>779</ID>
<type>AA_TOGGLE</type>
<position>39,-473</position>
<output>
<ID>OUT_0</ID>759 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>-76,-32</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>780</ID>
<type>AE_REGISTER8</type>
<position>63,-430</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>776 </input>
<input>
<ID>IN_2</ID>775 </input>
<input>
<ID>IN_3</ID>774 </input>
<input>
<ID>IN_4</ID>773 </input>
<input>
<ID>IN_5</ID>772 </input>
<input>
<ID>IN_6</ID>771 </input>
<input>
<ID>IN_7</ID>770 </input>
<input>
<ID>clock</ID>768 </input>
<input>
<ID>load</ID>769 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>-76,-44</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>781</ID>
<type>BB_CLOCK</type>
<position>62,-439</position>
<output>
<ID>CLK</ID>768 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>57,6.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>782</ID>
<type>AA_TOGGLE</type>
<position>62,-422</position>
<output>
<ID>OUT_0</ID>769 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>DE_TO</type>
<position>-76,-46</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>783</ID>
<type>AA_LABEL</type>
<position>68.5,-429.5</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>-76,-48</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>784</ID>
<type>AE_REGISTER8</type>
<position>40,-379</position>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>786 </input>
<input>
<ID>IN_2</ID>785 </input>
<input>
<ID>IN_3</ID>784 </input>
<input>
<ID>IN_4</ID>783 </input>
<input>
<ID>IN_5</ID>782 </input>
<input>
<ID>IN_6</ID>781 </input>
<input>
<ID>IN_7</ID>780 </input>
<input>
<ID>clock</ID>778 </input>
<input>
<ID>load</ID>779 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>-76,-42</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>785</ID>
<type>BB_CLOCK</type>
<position>39,-388</position>
<output>
<ID>CLK</ID>778 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>-32,21.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>786</ID>
<type>AA_TOGGLE</type>
<position>39,-371</position>
<output>
<ID>OUT_0</ID>779 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-32,19.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>787</ID>
<type>AA_LABEL</type>
<position>45.5,-378.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>-32,25.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>-39,30.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>-39,28.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>-39,26.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>-39,32.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>-80,-32</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>57,4.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-80,-34</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>57,2.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>-80,-36</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>57,0.5</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-80,-38</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>57,-11.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-80,-42</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>57,-13.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-80,-44</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>57,-15.5</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-80,-46</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>57,-17.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>-80,-48</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>65,-18</position>
<output>
<ID>A_greater_B</ID>26 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>103 </input>
<input>
<ID>IN_B_1</ID>104 </input>
<input>
<ID>IN_B_2</ID>105 </input>
<input>
<ID>IN_B_3</ID>106 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>-47,12</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>57,-29.5</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>-57,12</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>57,-31.5</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-67,12</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X3</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>57,-33.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>DA_FROM</type>
<position>-37,12</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID X0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>57,-35.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>-47,-23</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y1</lparam></gate>
<gate>
<ID>49</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>65,-36</position>
<output>
<ID>A_greater_B</ID>27 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>107 </input>
<input>
<ID>IN_B_1</ID>108 </input>
<input>
<ID>IN_B_2</ID>109 </input>
<input>
<ID>IN_B_3</ID>110 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>-57,-23</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y2</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>-67,-23</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y3</lparam></gate>
<gate>
<ID>52</ID>
<type>DA_FROM</type>
<position>-37,-23</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Y0</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_FULLADDER_4BIT</type>
<position>47,-13</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>97 </input>
<input>
<ID>IN_B_0</ID>115 </input>
<input>
<ID>IN_B_1</ID>75 </input>
<input>
<ID>IN_B_2</ID>74 </input>
<input>
<ID>IN_B_3</ID>73 </input>
<output>
<ID>OUT_0</ID>111 </output>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>65,0</position>
<output>
<ID>A_greater_B</ID>28 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>99 </input>
<input>
<ID>IN_B_1</ID>100 </input>
<input>
<ID>IN_B_2</ID>101 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-24,26</position>
<output>
<ID>A_greater_B</ID>1 </output>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>4 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_B_0</ID>6 </input>
<input>
<ID>IN_B_1</ID>7 </input>
<input>
<ID>IN_B_2</ID>8 </input>
<input>
<ID>IN_B_3</ID>9 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_REGISTER4</type>
<position>75,-18.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>clock</ID>30 </input>
<input>
<ID>load</ID>29 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>74,-9.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>CC_PULSE</type>
<position>-75,-52</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>CC_PULSE</type>
<position>74,-26.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-78.5,-52</position>
<gparam>LABEL_TEXT pulse</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>74,-28</position>
<gparam>LABEL_TEXT update</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>84,-17.5</position>
<gparam>LABEL_TEXT blinds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>-87.5,-34.5</position>
<gparam>LABEL_TEXT outside</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>-86.5,-44.5</position>
<gparam>LABEL_TEXT inside</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>-68,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>-61,-12</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>-64,1</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>-66,-5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>-58,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>-54,1</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_OR2</type>
<position>-56,-5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_DFF_LOW</type>
<position>-51,-12</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>-48,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW</type>
<position>-41,-12</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>-44,1</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR2</type>
<position>-46,-5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>-38,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>-31,-12</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>-34,1</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR2</type>
<position>-36,-5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_SMALL_INVERTER</type>
<position>-45,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>-55,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>-65,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-89,-25</position>
<gparam>LABEL_TEXT shift/load</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-84,-25</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND2</type>
<position>-68,-33</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_DFF_LOW</type>
<position>-61,-46</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>-64,-33</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_OR2</type>
<position>-66,-39</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>-58,-33</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>-54,-33</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>-56,-39</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_DFF_LOW</type>
<position>-51,-46</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND2</type>
<position>-48,-33</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW</type>
<position>-41,-46</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>-44,-33</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>-46,-39</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>-38,-33</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_DFF_LOW</type>
<position>-31,-46</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>82 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>-34,-33</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_OR2</type>
<position>-36,-39</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>-35,-28</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>-45,-28</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>-55,-28</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_SMALL_INVERTER</type>
<position>-65,-28</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>-18,2</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>-18,-4</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>-69,-28</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>-69,6</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_SMALL_INVERTER</type>
<position>-23,-5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>-18,-14</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>-18,-20</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_SMALL_INVERTER</type>
<position>-23,-15</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_DFF_LOW</type>
<position>-1,-3</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_DFF_LOW</type>
<position>7,-3</position>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_DFF_LOW</type>
<position>15,-3</position>
<input>
<ID>IN_0</ID>74 </input>
<output>
<ID>OUT_0</ID>75 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_DFF_LOW</type>
<position>23,-3</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>115 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>-9,-1</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_DFF_LOW</type>
<position>-1,-19</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>77 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_DFF_LOW</type>
<position>7.5,-19</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>78 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_DFF_LOW</type>
<position>15.5,-19</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-19</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_OR2</type>
<position>-9,-17</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>-26.5,-79.5</position>
<gparam>LABEL_TEXT loop activate-able</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>-80.5,-93</position>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-3.5,-97.5</position>
<gparam>LABEL_TEXT device 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-3.5,-110.5</position>
<gparam>LABEL_TEXT device 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_REGISTER4</type>
<position>-56.5,-104</position>
<output>
<ID>OUT_0</ID>121 </output>
<output>
<ID>OUT_1</ID>120 </output>
<output>
<ID>OUT_2</ID>119 </output>
<output>
<ID>OUT_3</ID>118 </output>
<input>
<ID>clear</ID>131 </input>
<input>
<ID>clock</ID>123 </input>
<input>
<ID>count_enable</ID>125 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND4</type>
<position>-47.5,-103.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>121 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>131</ID>
<type>BE_NOR2</type>
<position>-11.5,-92.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>BB_CLOCK</type>
<position>-63.5,-110</position>
<output>
<ID>CLK</ID>123 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 1</lparam></gate>
<gate>
<ID>133</ID>
<type>BE_NOR2</type>
<position>-11.5,-99.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>-5.5,-99.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>BE_NOR2</type>
<position>-65.5,-97</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>BE_NOR2</type>
<position>-65.5,-104</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>BE_NOR2</type>
<position>-37.5,-100</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>BE_NOR2</type>
<position>-37.5,-107</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_SMALL_INVERTER</type>
<position>-72.5,-105</position>
<input>
<ID>IN_0</ID>139 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>-86.5,-93</position>
<gparam>LABEL_TEXT occ. sensor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>-26.5,-82</position>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_OR2</type>
<position>-71.5,-96</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_OR2</type>
<position>-55.5,-113</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>-19.5,-94</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>-19.5,-98</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>-11.5,-105.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>BE_NOR2</type>
<position>-11.5,-112.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>-5.5,-112.5</position>
<input>
<ID>N_in0</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>-19.5,-107</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>-19.5,-111</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_SMALL_INVERTER</type>
<position>-24.5,-88</position>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_AND2</type>
<position>-79,-211</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>-86,-161.5</position>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-202.5</position>
<input>
<ID>IN_0</ID>401 </input>
<output>
<ID>OUT_0</ID>399 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-198.5</position>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>401 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>AE_SMALL_INVERTER</type>
<position>112.5,-215</position>
<input>
<ID>IN_0</ID>260 </input>
<output>
<ID>OUT_0</ID>402 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>-93,-161</position>
<gparam>LABEL_TEXT Change Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AE_SMALL_INVERTER</type>
<position>114.5,-298</position>
<input>
<ID>IN_0</ID>260 </input>
<output>
<ID>OUT_0</ID>403 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>50.5,-181.5</position>
<input>
<ID>N_in0</ID>140 </input>
<input>
<ID>N_in1</ID>202 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND4</type>
<position>46.5,-181.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>148 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>50.5,-189.5</position>
<input>
<ID>N_in0</ID>141 </input>
<input>
<ID>N_in1</ID>212 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND4</type>
<position>46.5,-189.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>50.5,-197.5</position>
<input>
<ID>N_in0</ID>142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND4</type>
<position>46.5,-197.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>148 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>50.5,-205.5</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_AND4</type>
<position>46.5,-205.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>50.5,-213.5</position>
<input>
<ID>N_in0</ID>144 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND4</type>
<position>46.5,-213.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>148 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>50.5,-221.5</position>
<input>
<ID>N_in0</ID>145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND4</type>
<position>46.5,-221.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>171</ID>
<type>GA_LED</type>
<position>50.5,-229.5</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND4</type>
<position>46.5,-229.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>148 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>50.5,-237.5</position>
<input>
<ID>N_in0</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND4</type>
<position>46.5,-237.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>153 </input>
<input>
<ID>IN_3</ID>152 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>-65,-229</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>259 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_SMALL_INVERTER</type>
<position>31.5,-170.5</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>177</ID>
<type>AE_SMALL_INVERTER</type>
<position>35,-170.5</position>
<input>
<ID>IN_0</ID>153 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_SMALL_INVERTER</type>
<position>38.5,-170.5</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_DFF_LOW</type>
<position>-53.5,-205</position>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>158 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>-51,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-214</position>
<input>
<ID>IN_0</ID>399 </input>
<output>
<ID>OUT_0</ID>269 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>-47,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR2</type>
<position>-49,-198</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AE_SMALL_INVERTER</type>
<position>-94,-218</position>
<input>
<ID>IN_0</ID>269 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR2</type>
<position>-71.5,-223.5</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_SMALL_INVERTER</type>
<position>-56.5,-188.5</position>
<input>
<ID>IN_0</ID>308 </input>
<output>
<ID>OUT_0</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AE_DFF_LOW</type>
<position>-44.5,-205</position>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>161 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>188</ID>
<type>AE_SMALL_INVERTER</type>
<position>-79.5,-231</position>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_AND2</type>
<position>-42,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>-38,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_OR2</type>
<position>-40,-198</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AE_DFF_LOW</type>
<position>-35.5,-205</position>
<input>
<ID>IN_0</ID>181 </input>
<output>
<ID>OUT_0</ID>164 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>193</ID>
<type>AA_AND2</type>
<position>-33,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_AND2</type>
<position>-29,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_OR2</type>
<position>-31,-198</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_DFF_LOW</type>
<position>-26,-205</position>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>167 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_AND2</type>
<position>-23.5,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>167 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>-19.5,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>189 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_OR2</type>
<position>-21.5,-198</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_DFF_LOW</type>
<position>-17,-205</position>
<input>
<ID>IN_0</ID>182 </input>
<output>
<ID>OUT_0</ID>170 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>-14.5,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND2</type>
<position>-10.5,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_OR2</type>
<position>-12.5,-198</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_DFF_LOW</type>
<position>-8,-205</position>
<input>
<ID>IN_0</ID>183 </input>
<output>
<ID>OUT_0</ID>173 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>-5.5,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>-1.5,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_OR2</type>
<position>-3.5,-198</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_DFF_LOW</type>
<position>1,-205</position>
<input>
<ID>IN_0</ID>184 </input>
<output>
<ID>OUT_0</ID>176 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND2</type>
<position>3.5,-192</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND2</type>
<position>7.5,-192</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_OR2</type>
<position>5.5,-198</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>174 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_DFF_LOW</type>
<position>10,-205</position>
<input>
<ID>IN_0</ID>185 </input>
<output>
<ID>OUT_0</ID>151 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_REGISTER8</type>
<position>-66.5,-182.5</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<input>
<ID>IN_2</ID>228 </input>
<input>
<ID>IN_3</ID>227 </input>
<input>
<ID>IN_4</ID>226 </input>
<input>
<ID>IN_5</ID>225 </input>
<input>
<ID>IN_6</ID>224 </input>
<input>
<ID>IN_7</ID>223 </input>
<output>
<ID>OUT_0</ID>177 </output>
<output>
<ID>OUT_1</ID>178 </output>
<output>
<ID>OUT_2</ID>191 </output>
<output>
<ID>OUT_3</ID>190 </output>
<output>
<ID>OUT_4</ID>189 </output>
<output>
<ID>OUT_5</ID>188 </output>
<output>
<ID>OUT_6</ID>187 </output>
<output>
<ID>OUT_7</ID>186 </output>
<input>
<ID>clock</ID>273 </input>
<input>
<ID>load</ID>231 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>214</ID>
<type>BB_CLOCK</type>
<position>-92.5,-229</position>
<output>
<ID>CLK</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>-77,-226.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_REGISTER4</type>
<position>-78.5,-218.5</position>
<output>
<ID>OUT_0</ID>232 </output>
<output>
<ID>OUT_3</ID>201 </output>
<input>
<ID>clear</ID>200 </input>
<input>
<ID>clock</ID>198 </input>
<input>
<ID>count_enable</ID>199 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-218.5</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_SMALL_INVERTER</type>
<position>-88.5,-223.5</position>
<input>
<ID>IN_0</ID>200 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND2</type>
<position>-83.5,-224.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AE_REGISTER8</type>
<position>113.5,-208</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>205 </input>
<input>
<ID>IN_3</ID>206 </input>
<input>
<ID>IN_4</ID>207 </input>
<input>
<ID>IN_5</ID>208 </input>
<input>
<ID>IN_6</ID>209 </input>
<input>
<ID>IN_7</ID>210 </input>
<output>
<ID>OUT_0</ID>381 </output>
<output>
<ID>OUT_1</ID>382 </output>
<output>
<ID>OUT_2</ID>383 </output>
<output>
<ID>OUT_3</ID>384 </output>
<output>
<ID>OUT_4</ID>385 </output>
<output>
<ID>OUT_5</ID>404 </output>
<output>
<ID>OUT_6</ID>387 </output>
<output>
<ID>OUT_7</ID>388 </output>
<input>
<ID>clock</ID>402 </input>
<input>
<ID>load</ID>211 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>221</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-234</position>
<input>
<ID>IN_0</ID>202 </input>
<output>
<ID>OUT_0</ID>203 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>222</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-225.5</position>
<input>
<ID>IN_0</ID>203 </input>
<output>
<ID>OUT_0</ID>204 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-217</position>
<input>
<ID>IN_0</ID>204 </input>
<output>
<ID>OUT_0</ID>205 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-209</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUT_0</ID>206 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-201.5</position>
<input>
<ID>IN_0</ID>206 </input>
<output>
<ID>OUT_0</ID>207 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>226</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-194</position>
<input>
<ID>IN_0</ID>207 </input>
<output>
<ID>OUT_0</ID>208 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-186.5</position>
<input>
<ID>IN_0</ID>208 </input>
<output>
<ID>OUT_0</ID>209 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_DFF_LOW</type>
<position>86.5,-179</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>210 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_TOGGLE</type>
<position>112.5,-200</position>
<output>
<ID>OUT_0</ID>211 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_REGISTER8</type>
<position>115.5,-291</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<input>
<ID>IN_2</ID>215 </input>
<input>
<ID>IN_3</ID>216 </input>
<input>
<ID>IN_4</ID>217 </input>
<input>
<ID>IN_5</ID>218 </input>
<input>
<ID>IN_6</ID>219 </input>
<input>
<ID>IN_7</ID>220 </input>
<output>
<ID>OUT_0</ID>389 </output>
<output>
<ID>OUT_1</ID>390 </output>
<output>
<ID>OUT_2</ID>391 </output>
<output>
<ID>OUT_3</ID>392 </output>
<output>
<ID>OUT_4</ID>393 </output>
<output>
<ID>OUT_5</ID>394 </output>
<output>
<ID>OUT_6</ID>395 </output>
<output>
<ID>OUT_7</ID>380 </output>
<input>
<ID>clock</ID>403 </input>
<input>
<ID>load</ID>222 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 128</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>231</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-317</position>
<input>
<ID>IN_0</ID>212 </input>
<output>
<ID>OUT_0</ID>213 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-308.5</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>214 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>233</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-300</position>
<input>
<ID>IN_0</ID>214 </input>
<output>
<ID>OUT_0</ID>215 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>234</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-292</position>
<input>
<ID>IN_0</ID>215 </input>
<output>
<ID>OUT_0</ID>216 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>235</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-284.5</position>
<input>
<ID>IN_0</ID>216 </input>
<output>
<ID>OUT_0</ID>217 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>236</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-277</position>
<input>
<ID>IN_0</ID>217 </input>
<output>
<ID>OUT_0</ID>218 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>237</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-269.5</position>
<input>
<ID>IN_0</ID>218 </input>
<output>
<ID>OUT_0</ID>219 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_DFF_LOW</type>
<position>88.5,-262</position>
<input>
<ID>IN_0</ID>219 </input>
<output>
<ID>OUT_0</ID>220 </output>
<input>
<ID>clock</ID>260 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>-74.5,-203</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_TOGGLE</type>
<position>114.5,-283</position>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-176.5</position>
<output>
<ID>OUT_0</ID>223 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-178.5</position>
<output>
<ID>OUT_0</ID>224 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-180.5</position>
<output>
<ID>OUT_0</ID>225 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-182.5</position>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-184.5</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-186.5</position>
<output>
<ID>OUT_0</ID>228 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-188.5</position>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>-85.5,-190.5</position>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>-67.5,-174.5</position>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>-91.5,-183.5</position>
<gparam>LABEL_TEXT New Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND2</type>
<position>-57,-228</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>AE_OR2</type>
<position>-86,-196.5</position>
<input>
<ID>IN_0</ID>407 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>-57,-236</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>407 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>-47.5,-222.5</position>
<input>
<ID>IN_0</ID>407 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>271 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AE_SMALL_INVERTER</type>
<position>-31,-219</position>
<input>
<ID>IN_0</ID>268 </input>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>256</ID>
<type>AI_MUX_8x1</type>
<position>233.5,-262.5</position>
<input>
<ID>IN_0</ID>406 </input>
<input>
<ID>IN_1</ID>405 </input>
<output>
<ID>OUT</ID>234 </output>
<input>
<ID>SEL_0</ID>152 </input>
<input>
<ID>SEL_1</ID>153 </input>
<input>
<ID>SEL_2</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_MUX_2x1</type>
<position>358,-260</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>367 </output>
<input>
<ID>SEL_0</ID>407 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>281.5,-275.5</position>
<gparam>LABEL_TEXT Default</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>310,-256</position>
<gparam>LABEL_TEXT Custom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>395.5,-249.5</position>
<gparam>LABEL_TEXT Light</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AE_DFF_LOW</type>
<position>152.5,-290.5</position>
<input>
<ID>IN_0</ID>389 </input>
<output>
<ID>OUT_0</ID>240 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>155,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_AND2</type>
<position>159,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>390 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_OR2</type>
<position>157,-283.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>-30,-222.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AE_SMALL_INVERTER</type>
<position>-36.5,-222.5</position>
<input>
<ID>IN_0</ID>271 </input>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_DFF_LOW</type>
<position>161.5,-290.5</position>
<input>
<ID>IN_0</ID>261 </input>
<output>
<ID>OUT_0</ID>243 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_AND2</type>
<position>164,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>241 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_AND2</type>
<position>168,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>391 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_OR2</type>
<position>166,-283.5</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AE_DFF_LOW</type>
<position>170.5,-290.5</position>
<input>
<ID>IN_0</ID>263 </input>
<output>
<ID>OUT_0</ID>246 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_AND2</type>
<position>173,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_AND2</type>
<position>177,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>392 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_OR2</type>
<position>175,-283.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>AE_DFF_LOW</type>
<position>180,-290.5</position>
<input>
<ID>IN_0</ID>262 </input>
<output>
<ID>OUT_0</ID>249 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>182.5,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>186.5,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>393 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AE_OR2</type>
<position>184.5,-283.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>264 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AE_DFF_LOW</type>
<position>189,-290.5</position>
<input>
<ID>IN_0</ID>264 </input>
<output>
<ID>OUT_0</ID>252 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>191.5,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>195.5,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>394 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_OR2</type>
<position>193.5,-283.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>265 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>AE_DFF_LOW</type>
<position>198,-290.5</position>
<input>
<ID>IN_0</ID>265 </input>
<output>
<ID>OUT_0</ID>255 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_AND2</type>
<position>200.5,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>AA_AND2</type>
<position>204.5,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>395 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_OR2</type>
<position>202.5,-283.5</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>AE_DFF_LOW</type>
<position>207,-290.5</position>
<input>
<ID>IN_0</ID>266 </input>
<output>
<ID>OUT_0</ID>258 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND2</type>
<position>209.5,-277.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>256 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_AND2</type>
<position>213.5,-277.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>380 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_OR2</type>
<position>211.5,-283.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_DFF_LOW</type>
<position>216,-290.5</position>
<input>
<ID>IN_0</ID>267 </input>
<output>
<ID>OUT_0</ID>405 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>292</ID>
<type>BB_CLOCK</type>
<position>-70.5,-191.5</position>
<output>
<ID>CLK</ID>273 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>293</ID>
<type>AA_AND2</type>
<position>-63.5,-194.5</position>
<input>
<ID>IN_0</ID>308 </input>
<input>
<ID>IN_1</ID>308 </input>
<output>
<ID>OUT</ID>272 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_DFF_LOW</type>
<position>151,-231</position>
<input>
<ID>IN_0</ID>381 </input>
<output>
<ID>OUT_0</ID>278 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND2</type>
<position>153.5,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>278 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>239.5,-305.5</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>312 </input>
<output>
<ID>OUT</ID>310 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_AND2</type>
<position>157.5,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>382 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>AE_OR2</type>
<position>155.5,-224</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>AE_SMALL_INVERTER</type>
<position>229,-293.5</position>
<input>
<ID>IN_0</ID>319 </input>
<output>
<ID>OUT_0</ID>317 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_SMALL_INVERTER</type>
<position>229,-289.5</position>
<input>
<ID>IN_0</ID>379 </input>
<output>
<ID>OUT_0</ID>319 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND2</type>
<position>254.5,-321</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>314 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_DFF_LOW</type>
<position>160,-231</position>
<input>
<ID>IN_0</ID>299 </input>
<output>
<ID>OUT_0</ID>281 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_SMALL_INVERTER</type>
<position>224.5,-308.5</position>
<input>
<ID>IN_0</ID>317 </input>
<output>
<ID>OUT_0</ID>315 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>162.5,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>281 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>166.5,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>383 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_OR2</type>
<position>164.5,-224</position>
<input>
<ID>IN_0</ID>280 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_DFF_LOW</type>
<position>169,-231</position>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>284 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND2</type>
<position>171.5,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_AND2</type>
<position>175.5,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>384 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>310</ID>
<type>AE_OR2</type>
<position>173.5,-224</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>282 </input>
<output>
<ID>OUT</ID>300 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-231</position>
<input>
<ID>IN_0</ID>300 </input>
<output>
<ID>OUT_0</ID>287 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_AND2</type>
<position>181,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>185,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>286 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>AE_OR2</type>
<position>183,-224</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>285 </input>
<output>
<ID>OUT</ID>302 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>AE_DFF_LOW</type>
<position>187.5,-231</position>
<input>
<ID>IN_0</ID>302 </input>
<output>
<ID>OUT_0</ID>290 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_AND2</type>
<position>190,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_AND2</type>
<position>194,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>404 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AE_OR2</type>
<position>192,-224</position>
<input>
<ID>IN_0</ID>289 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>303 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_DFF_LOW</type>
<position>196.5,-231</position>
<input>
<ID>IN_0</ID>303 </input>
<output>
<ID>OUT_0</ID>293 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>199,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>293 </input>
<output>
<ID>OUT</ID>291 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_AND2</type>
<position>203,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>387 </input>
<output>
<ID>OUT</ID>292 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>AE_OR2</type>
<position>201,-224</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>291 </input>
<output>
<ID>OUT</ID>304 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_DFF_LOW</type>
<position>205.5,-231</position>
<input>
<ID>IN_0</ID>304 </input>
<output>
<ID>OUT_0</ID>296 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_AND2</type>
<position>208,-218</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>294 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND2</type>
<position>212,-218</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>295 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_OR2</type>
<position>210,-224</position>
<input>
<ID>IN_0</ID>295 </input>
<input>
<ID>IN_1</ID>294 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AE_DFF_LOW</type>
<position>214.5,-231</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>406 </output>
<input>
<ID>clock</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_SMALL_INVERTER</type>
<position>224.5,-312.5</position>
<input>
<ID>IN_0</ID>315 </input>
<output>
<ID>OUT_0</ID>298 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>329</ID>
<type>AE_OR2</type>
<position>247,-318</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>306 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AE_SMALL_INVERTER</type>
<position>239,-325.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>BB_CLOCK</type>
<position>226,-323.5</position>
<output>
<ID>CLK</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_AND2</type>
<position>241.5,-321</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>276 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_REGISTER4</type>
<position>240,-313</position>
<output>
<ID>OUT_0</ID>312 </output>
<output>
<ID>OUT_3</ID>311 </output>
<input>
<ID>clear</ID>310 </input>
<input>
<ID>clock</ID>307 </input>
<input>
<ID>count_enable</ID>309 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>233,-313</position>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_SMALL_INVERTER</type>
<position>230,-318</position>
<input>
<ID>IN_0</ID>310 </input>
<output>
<ID>OUT_0</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_AND2</type>
<position>235,-319</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_DFF_LOW</type>
<position>266,-307.5</position>
<input>
<ID>IN_0</ID>343 </input>
<output>
<ID>OUT_0</ID>324 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>268.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_AND2</type>
<position>272.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>397 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AE_OR2</type>
<position>270.5,-300.5</position>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>344 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AA_AND2</type>
<position>254,-297.5</position>
<input>
<ID>IN_0</ID>316 </input>
<input>
<ID>IN_1</ID>316 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_DFF_LOW</type>
<position>275,-307.5</position>
<input>
<ID>IN_0</ID>344 </input>
<output>
<ID>OUT_0</ID>327 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>277.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_AND2</type>
<position>281.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>356 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AE_OR2</type>
<position>279.5,-300.5</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>346 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_DFF_LOW</type>
<position>284,-307.5</position>
<input>
<ID>IN_0</ID>346 </input>
<output>
<ID>OUT_0</ID>330 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>347</ID>
<type>AA_AND2</type>
<position>286.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>328 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_AND2</type>
<position>290.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>329 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AE_OR2</type>
<position>288.5,-300.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_DFF_LOW</type>
<position>293.5,-307.5</position>
<input>
<ID>IN_0</ID>345 </input>
<output>
<ID>OUT_0</ID>333 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND2</type>
<position>295.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>331 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND2</type>
<position>299.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>354 </input>
<output>
<ID>OUT</ID>332 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_OR2</type>
<position>297.5,-300.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<output>
<ID>OUT</ID>347 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AE_DFF_LOW</type>
<position>302,-307.5</position>
<input>
<ID>IN_0</ID>347 </input>
<output>
<ID>OUT_0</ID>336 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>304.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>336 </input>
<output>
<ID>OUT</ID>334 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_AND2</type>
<position>308.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>353 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AE_OR2</type>
<position>306.5,-300.5</position>
<input>
<ID>IN_0</ID>335 </input>
<input>
<ID>IN_1</ID>334 </input>
<output>
<ID>OUT</ID>348 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AE_DFF_LOW</type>
<position>311,-307.5</position>
<input>
<ID>IN_0</ID>348 </input>
<output>
<ID>OUT_0</ID>339 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>313.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>339 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>317.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AE_OR2</type>
<position>315.5,-300.5</position>
<input>
<ID>IN_0</ID>338 </input>
<input>
<ID>IN_1</ID>337 </input>
<output>
<ID>OUT</ID>349 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AE_DFF_LOW</type>
<position>320,-307.5</position>
<input>
<ID>IN_0</ID>349 </input>
<output>
<ID>OUT_0</ID>342 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>322.5,-294.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>342 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AA_AND2</type>
<position>326.5,-294.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_OR2</type>
<position>324.5,-300.5</position>
<input>
<ID>IN_0</ID>341 </input>
<input>
<ID>IN_1</ID>340 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_DFF_LOW</type>
<position>329,-307.5</position>
<input>
<ID>IN_0</ID>350 </input>
<output>
<ID>OUT_0</ID>377 </output>
<input>
<ID>clock</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>367</ID>
<type>AE_SMALL_INVERTER</type>
<position>230,-299.5</position>
<input>
<ID>IN_0</ID>317 </input>
<output>
<ID>OUT_0</ID>318 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_REGISTER8</type>
<position>253,-285</position>
<input>
<ID>IN_0</ID>358 </input>
<input>
<ID>IN_1</ID>359 </input>
<input>
<ID>IN_2</ID>360 </input>
<input>
<ID>IN_3</ID>361 </input>
<input>
<ID>IN_4</ID>362 </input>
<input>
<ID>IN_5</ID>364 </input>
<input>
<ID>IN_6</ID>363 </input>
<input>
<ID>IN_7</ID>365 </input>
<output>
<ID>OUT_0</ID>343 </output>
<output>
<ID>OUT_1</ID>397 </output>
<output>
<ID>OUT_2</ID>356 </output>
<output>
<ID>OUT_3</ID>355 </output>
<output>
<ID>OUT_4</ID>354 </output>
<output>
<ID>OUT_5</ID>353 </output>
<output>
<ID>OUT_6</ID>352 </output>
<output>
<ID>OUT_7</ID>351 </output>
<input>
<ID>clock</ID>357 </input>
<input>
<ID>load</ID>366 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 135</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_TOGGLE</type>
<position>252,-292</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_TOGGLE</type>
<position>252,-277</position>
<output>
<ID>OUT_0</ID>366 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_TOGGLE</type>
<position>241,-277.5</position>
<output>
<ID>OUT_0</ID>365 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_TOGGLE</type>
<position>241,-279.5</position>
<output>
<ID>OUT_0</ID>363 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>373</ID>
<type>AA_TOGGLE</type>
<position>241,-281.5</position>
<output>
<ID>OUT_0</ID>364 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_TOGGLE</type>
<position>241,-283.5</position>
<output>
<ID>OUT_0</ID>362 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_TOGGLE</type>
<position>241,-285.5</position>
<output>
<ID>OUT_0</ID>361 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>376</ID>
<type>AA_TOGGLE</type>
<position>241,-287.5</position>
<output>
<ID>OUT_0</ID>360 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_TOGGLE</type>
<position>241,-289.5</position>
<output>
<ID>OUT_0</ID>359 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_TOGGLE</type>
<position>241,-291.5</position>
<output>
<ID>OUT_0</ID>358 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_REGISTER8</type>
<position>388,-251</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>369 </input>
<input>
<ID>IN_2</ID>370 </input>
<input>
<ID>IN_3</ID>371 </input>
<input>
<ID>IN_4</ID>372 </input>
<input>
<ID>IN_5</ID>373 </input>
<input>
<ID>IN_6</ID>374 </input>
<input>
<ID>IN_7</ID>375 </input>
<input>
<ID>clock</ID>398 </input>
<input>
<ID>load</ID>376 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 128</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_DFF_LOW</type>
<position>374,-279</position>
<input>
<ID>IN_0</ID>367 </input>
<output>
<ID>OUT_0</ID>368 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>381</ID>
<type>AE_DFF_LOW</type>
<position>374,-271</position>
<input>
<ID>IN_0</ID>368 </input>
<output>
<ID>OUT_0</ID>369 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>382</ID>
<type>AE_DFF_LOW</type>
<position>374,-263</position>
<input>
<ID>IN_0</ID>369 </input>
<output>
<ID>OUT_0</ID>370 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_DFF_LOW</type>
<position>374,-255</position>
<input>
<ID>IN_0</ID>370 </input>
<output>
<ID>OUT_0</ID>371 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>384</ID>
<type>AE_DFF_LOW</type>
<position>374,-247</position>
<input>
<ID>IN_0</ID>371 </input>
<output>
<ID>OUT_0</ID>372 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>385</ID>
<type>AE_DFF_LOW</type>
<position>374,-239</position>
<input>
<ID>IN_0</ID>372 </input>
<output>
<ID>OUT_0</ID>373 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>386</ID>
<type>AE_DFF_LOW</type>
<position>374,-231</position>
<input>
<ID>IN_0</ID>373 </input>
<output>
<ID>OUT_0</ID>374 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>387</ID>
<type>AE_DFF_LOW</type>
<position>374,-223</position>
<input>
<ID>IN_0</ID>374 </input>
<output>
<ID>OUT_0</ID>375 </output>
<input>
<ID>clock</ID>396 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_TOGGLE</type>
<position>387,-243</position>
<output>
<ID>OUT_0</ID>376 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>389</ID>
<type>AE_SMALL_INVERTER</type>
<position>387,-258</position>
<input>
<ID>IN_0</ID>396 </input>
<output>
<ID>OUT_0</ID>398 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_AND2</type>
<position>235,-298.5</position>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>AE_SMALL_INVERTER</type>
<position>249,-298.5</position>
<input>
<ID>IN_0</ID>313 </input>
<output>
<ID>OUT_0</ID>316 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>392</ID>
<type>AE_SMALL_INVERTER</type>
<position>260.5,-290.5</position>
<input>
<ID>IN_0</ID>316 </input>
<output>
<ID>OUT_0</ID>378 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>393</ID>
<type>AA_TOGGLE</type>
<position>-86,-158.5</position>
<output>
<ID>OUT_0</ID>407 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_TOGGLE</type>
<position>-86,-164.5</position>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_TOGGLE</type>
<position>-86,-166.5</position>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_TOGGLE</type>
<position>-86,-168.5</position>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_LABEL</type>
<position>-89.5,-158.5</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>398</ID>
<type>AA_LABEL</type>
<position>-92.5,-166.5</position>
<gparam>LABEL_TEXT Notif Index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>399</ID>
<type>AE_SMALL_INVERTER</type>
<position>235,-287.5</position>
<input>
<ID>IN_0</ID>407 </input>
<output>
<ID>OUT_0</ID>379 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>368.5,-304.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>320 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>401</ID>
<type>AE_SMALL_INVERTER</type>
<position>-88.5,-205</position>
<input>
<ID>IN_0</ID>399 </input>
<output>
<ID>OUT_0</ID>400 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>402</ID>
<type>AA_AND2</type>
<position>-83.5,-204</position>
<input>
<ID>IN_0</ID>399 </input>
<input>
<ID>IN_1</ID>400 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AE_SMALL_INVERTER</type>
<position>-69.5,-195.5</position>
<input>
<ID>IN_0</ID>233 </input>
<output>
<ID>OUT_0</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_TOGGLE</type>
<position>-73,84.5</position>
<output>
<ID>OUT_0</ID>423 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_TOGGLE</type>
<position>-73,80.5</position>
<output>
<ID>OUT_0</ID>408 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_TOGGLE</type>
<position>-73,76.5</position>
<output>
<ID>OUT_0</ID>409 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>407</ID>
<type>AE_OR2</type>
<position>-66,78.5</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>-58,77.5</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>413 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_TOGGLE</type>
<position>-73,70.5</position>
<output>
<ID>OUT_0</ID>412 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_OR2</type>
<position>-50,83.5</position>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>411 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_LABEL</type>
<position>-78,84.5</position>
<gparam>LABEL_TEXT mag. lock</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>412</ID>
<type>AA_LABEL</type>
<position>-79.5,80.5</position>
<gparam>LABEL_TEXT sound sensor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>AA_LABEL</type>
<position>-78.5,76.5</position>
<gparam>LABEL_TEXT occ. sensor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AA_LABEL</type>
<position>-76,70.5</position>
<gparam>LABEL_TEXT GPS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>AA_INVERTER</type>
<position>-66,70.5</position>
<input>
<ID>IN_0</ID>412 </input>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>416</ID>
<type>BE_NOR2</type>
<position>-42,82.5</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>418 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>BE_NOR2</type>
<position>-42,75.5</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>-76.5,61.5</position>
<gparam>LABEL_TEXT reset</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>CC_PULSE</type>
<position>-73,61.5</position>
<output>
<ID>OUT_0</ID>417 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>GA_LED</type>
<position>-33,75.5</position>
<input>
<ID>N_in0</ID>418 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>421</ID>
<type>AA_LABEL</type>
<position>-21.5,75.5</position>
<gparam>LABEL_TEXT alarm, police, video, notify</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>GA_LED</type>
<position>-19,60.5</position>
<input>
<ID>N_in0</ID>422 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>BE_NOR2</type>
<position>-26,67.5</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>422 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>424</ID>
<type>BE_NOR2</type>
<position>-26,60.5</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>CC_PULSE</type>
<position>-49,63.5</position>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AE_OR2</type>
<position>-42,62.5</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_LABEL</type>
<position>-53.5,63.5</position>
<gparam>LABEL_TEXT hang up</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_LABEL</type>
<position>-13,60.5</position>
<gparam>LABEL_TEXT conversation</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_AND2</type>
<position>-34,68.5</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>CC_PULSE</type>
<position>-49,67.5</position>
<output>
<ID>OUT_0</ID>419 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_LABEL</type>
<position>-51.5,67.5</position>
<gparam>LABEL_TEXT call</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>606</ID>
<type>AA_TOGGLE</type>
<position>-52,-407</position>
<output>
<ID>OUT_0</ID>804 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_LABEL</type>
<position>-56,-407</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>608</ID>
<type>BE_JKFF_LOW</type>
<position>-53,-389</position>
<input>
<ID>J</ID>594 </input>
<input>
<ID>K</ID>594 </input>
<output>
<ID>Q</ID>751 </output>
<input>
<ID>clear</ID>804 </input>
<input>
<ID>clock</ID>595 </input>
<output>
<ID>nQ</ID>597 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>609</ID>
<type>BE_JKFF_LOW</type>
<position>-22,-389</position>
<input>
<ID>J</ID>600 </input>
<input>
<ID>K</ID>600 </input>
<output>
<ID>Q</ID>695 </output>
<input>
<ID>clear</ID>804 </input>
<input>
<ID>clock</ID>595 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_TOGGLE</type>
<position>-61,-387</position>
<output>
<ID>OUT_0</ID>594 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>611</ID>
<type>AA_LABEL</type>
<position>-65,-386.5</position>
<gparam>LABEL_TEXT Logic1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>612</ID>
<type>AA_AND2</type>
<position>-38,-387</position>
<input>
<ID>IN_0</ID>604 </input>
<input>
<ID>IN_1</ID>751 </input>
<output>
<ID>OUT</ID>598 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_AND2</type>
<position>-38,-391</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>596 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>614</ID>
<type>AE_SMALL_INVERTER</type>
<position>-46,-392</position>
<input>
<ID>IN_0</ID>604 </input>
<output>
<ID>OUT_0</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>615</ID>
<type>AE_OR2</type>
<position>-30,-389</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>599 </input>
<output>
<ID>OUT</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_LABEL</type>
<position>-29.5,-363.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>617</ID>
<type>AA_LABEL</type>
<position>-25,-412.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>618</ID>
<type>AA_TOGGLE</type>
<position>-52,-403</position>
<output>
<ID>OUT_0</ID>601 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>619</ID>
<type>AA_TOGGLE</type>
<position>-52,-401</position>
<output>
<ID>OUT_0</ID>604 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>621</ID>
<type>AA_LABEL</type>
<position>-56,-403</position>
<gparam>LABEL_TEXT Update</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>622</ID>
<type>AA_LABEL</type>
<position>-60.5,-401</position>
<gparam>LABEL_TEXT Increase/Decrease</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>623</ID>
<type>AE_SMALL_INVERTER</type>
<position>-17,-405</position>
<input>
<ID>IN_0</ID>602 </input>
<output>
<ID>OUT_0</ID>603 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>624</ID>
<type>AA_LABEL</type>
<position>-26,-403</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>625</ID>
<type>AA_TOGGLE</type>
<position>-22,-403</position>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>626</ID>
<type>AE_REGISTER8</type>
<position>-17,-413</position>
<output>
<ID>OUT_0</ID>612 </output>
<output>
<ID>OUT_1</ID>611 </output>
<output>
<ID>OUT_2</ID>610 </output>
<output>
<ID>OUT_3</ID>609 </output>
<output>
<ID>OUT_4</ID>608 </output>
<output>
<ID>OUT_5</ID>607 </output>
<output>
<ID>OUT_6</ID>606 </output>
<output>
<ID>OUT_7</ID>605 </output>
<output>
<ID>carry_out</ID>595 </output>
<input>
<ID>clear</ID>804 </input>
<input>
<ID>clock</ID>601 </input>
<input>
<ID>count_enable</ID>603 </input>
<input>
<ID>count_up</ID>604 </input>
<input>
<ID>load</ID>602 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>627</ID>
<type>AA_LABEL</type>
<position>-4.5,-359</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>639</ID>
<type>AA_LABEL</type>
<position>45.5,-480.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>640</ID>
<type>AE_OR2</type>
<position>47,-415.5</position>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>795 </input>
<output>
<ID>OUT</ID>777 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>AE_OR2</type>
<position>47,-419.5</position>
<input>
<ID>IN_0</ID>797 </input>
<input>
<ID>IN_1</ID>794 </input>
<output>
<ID>OUT</ID>776 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>642</ID>
<type>AE_OR2</type>
<position>47,-423.5</position>
<input>
<ID>IN_0</ID>798 </input>
<input>
<ID>IN_1</ID>793 </input>
<output>
<ID>OUT</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>643</ID>
<type>AE_OR2</type>
<position>47,-427.5</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>792 </input>
<output>
<ID>OUT</ID>774 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>AE_OR2</type>
<position>47,-431.5</position>
<input>
<ID>IN_0</ID>800 </input>
<input>
<ID>IN_1</ID>791 </input>
<output>
<ID>OUT</ID>773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>645</ID>
<type>AE_OR2</type>
<position>47,-435.5</position>
<input>
<ID>IN_0</ID>801 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>646</ID>
<type>AE_OR2</type>
<position>47,-439.5</position>
<input>
<ID>IN_0</ID>802 </input>
<input>
<ID>IN_1</ID>789 </input>
<output>
<ID>OUT</ID>771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>647</ID>
<type>AE_OR2</type>
<position>47,-443.5</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>788 </input>
<output>
<ID>OUT</ID>770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_AND2</type>
<position>24,-364.5</position>
<input>
<ID>IN_0</ID>637 </input>
<input>
<ID>IN_1</ID>638 </input>
<output>
<ID>OUT</ID>787 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-363.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>637 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>651</ID>
<type>AA_AND2</type>
<position>24,-368.5</position>
<input>
<ID>IN_0</ID>668 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>786 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_AND2</type>
<position>24,-372.5</position>
<input>
<ID>IN_0</ID>667 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>785 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>653</ID>
<type>AA_AND2</type>
<position>24,-376.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>784 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>654</ID>
<type>AA_AND2</type>
<position>24,-380.5</position>
<input>
<ID>IN_0</ID>665 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>655</ID>
<type>AA_AND2</type>
<position>24,-384.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>644 </input>
<output>
<ID>OUT</ID>782 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>AA_AND2</type>
<position>24,-388.5</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_AND2</type>
<position>24,-392.5</position>
<input>
<ID>IN_0</ID>662 </input>
<input>
<ID>IN_1</ID>646 </input>
<output>
<ID>OUT</ID>780 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>666</ID>
<type>AA_AND2</type>
<position>24,-398.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>638 </input>
<output>
<ID>OUT</ID>796 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_AND2</type>
<position>24,-402.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>797 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>668</ID>
<type>AA_AND2</type>
<position>24,-406.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>798 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>669</ID>
<type>AA_AND2</type>
<position>24,-410.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>799 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>AA_AND2</type>
<position>24,-414.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>800 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>671</ID>
<type>AA_AND2</type>
<position>24,-418.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>644 </input>
<output>
<ID>OUT</ID>801 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>672</ID>
<type>AA_AND2</type>
<position>24,-422.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>802 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>673</ID>
<type>AA_AND2</type>
<position>24,-426.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>646 </input>
<output>
<ID>OUT</ID>803 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>681</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-367.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>682</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-371.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>667 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>683</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-375.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>666 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>684</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-379.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>665 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>685</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-383.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>664 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>686</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-387.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>663 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-391.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>662 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_AND2</type>
<position>24,-432.5</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-431.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>669 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>691</ID>
<type>AA_AND2</type>
<position>24,-436.5</position>
<input>
<ID>IN_0</ID>701 </input>
<input>
<ID>IN_1</ID>672 </input>
<output>
<ID>OUT</ID>794 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>AA_AND2</type>
<position>24,-440.5</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>673 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>693</ID>
<type>AA_AND2</type>
<position>24,-444.5</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>674 </input>
<output>
<ID>OUT</ID>792 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>694</ID>
<type>AA_AND2</type>
<position>24,-448.5</position>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>791 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>AA_AND2</type>
<position>24,-452.5</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>676 </input>
<output>
<ID>OUT</ID>790 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>696</ID>
<type>AA_AND2</type>
<position>24,-456.5</position>
<input>
<ID>IN_0</ID>696 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>789 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_AND2</type>
<position>24,-460.5</position>
<input>
<ID>IN_0</ID>694 </input>
<input>
<ID>IN_1</ID>678 </input>
<output>
<ID>OUT</ID>788 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>706</ID>
<type>AA_AND2</type>
<position>24,-466.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>707</ID>
<type>AA_AND2</type>
<position>24,-470.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>672 </input>
<output>
<ID>OUT</ID>766 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>708</ID>
<type>AA_AND2</type>
<position>24,-474.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>673 </input>
<output>
<ID>OUT</ID>765 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>AA_AND2</type>
<position>24,-478.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>674 </input>
<output>
<ID>OUT</ID>764 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_AND2</type>
<position>24,-482.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>763 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>711</ID>
<type>AA_AND2</type>
<position>24,-486.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>676 </input>
<output>
<ID>OUT</ID>762 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>712</ID>
<type>AA_AND2</type>
<position>24,-490.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>713</ID>
<type>AA_AND2</type>
<position>24,-494.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>678 </input>
<output>
<ID>OUT</ID>760 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>721</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-435.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>701 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>722</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-439.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>723</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-443.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>699 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>724</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-447.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>725</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-451.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-455.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>696 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-459.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>694 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>744</ID>
<type>AA_LABEL</type>
<position>3,-361.5</position>
<gparam>LABEL_TEXT ~D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>745</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-366.5</position>
<input>
<ID>IN_0</ID>612 </input>
<output>
<ID>OUT_0</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>746</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-370.5</position>
<input>
<ID>IN_0</ID>611 </input>
<output>
<ID>OUT_0</ID>743 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>747</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-374.5</position>
<input>
<ID>IN_0</ID>610 </input>
<output>
<ID>OUT_0</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>748</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-378.5</position>
<input>
<ID>IN_0</ID>609 </input>
<output>
<ID>OUT_0</ID>745 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>749</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-382.5</position>
<input>
<ID>IN_0</ID>608 </input>
<output>
<ID>OUT_0</ID>746 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>750</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-386.5</position>
<input>
<ID>IN_0</ID>607 </input>
<output>
<ID>OUT_0</ID>747 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-390.5</position>
<input>
<ID>IN_0</ID>606 </input>
<output>
<ID>OUT_0</ID>748 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1,-394.5</position>
<input>
<ID>IN_0</ID>605 </input>
<output>
<ID>OUT_0</ID>749 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>753</ID>
<type>AE_OR2</type>
<position>4,-365.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>742 </input>
<output>
<ID>OUT</ID>638 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>754</ID>
<type>AE_OR2</type>
<position>4,-369.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>743 </input>
<output>
<ID>OUT</ID>640 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_OR2</type>
<position>4,-373.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>744 </input>
<output>
<ID>OUT</ID>641 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>756</ID>
<type>AE_OR2</type>
<position>4,-377.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>745 </input>
<output>
<ID>OUT</ID>642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>757</ID>
<type>AE_OR2</type>
<position>4,-381.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>746 </input>
<output>
<ID>OUT</ID>643 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>AE_OR2</type>
<position>4,-385.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>747 </input>
<output>
<ID>OUT</ID>644 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>759</ID>
<type>AE_OR2</type>
<position>4,-389.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>748 </input>
<output>
<ID>OUT</ID>645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>760</ID>
<type>AE_OR2</type>
<position>4,-393.5</position>
<input>
<ID>IN_0</ID>750 </input>
<input>
<ID>IN_1</ID>749 </input>
<output>
<ID>OUT</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AE_SMALL_INVERTER</type>
<position>-15,-364.5</position>
<input>
<ID>IN_0</ID>751 </input>
<output>
<ID>OUT_0</ID>750 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>762</ID>
<type>AA_LABEL</type>
<position>4,-429</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>763</ID>
<type>AE_OR2</type>
<position>4,-433.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>612 </input>
<output>
<ID>OUT</ID>670 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>764</ID>
<type>AE_OR2</type>
<position>4,-437.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>611 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>765</ID>
<type>AE_OR2</type>
<position>4,-441.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>610 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>AE_OR2</type>
<position>4,-445.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>609 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>767</ID>
<type>AE_OR2</type>
<position>4,-449.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>608 </input>
<output>
<ID>OUT</ID>675 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>768</ID>
<type>AE_OR2</type>
<position>4,-453.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>676 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>769</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>62,-424,62,-424</points>
<connection>
<GID>780</GID>
<name>load</name></connection>
<connection>
<GID>782</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-443.5,51,-426</points>
<intersection>-443.5 2</intersection>
<intersection>-426 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-426,59,-426</points>
<connection>
<GID>780</GID>
<name>IN_7</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-443.5,51,-443.5</points>
<connection>
<GID>647</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-21,-26,18</points>
<connection>
<GID>55</GID>
<name>A_greater_B</name></connection>
<intersection>-21 8</intersection>
<intersection>-15 10</intersection>
<intersection>-5 9</intersection>
<intersection>1 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-26,1,-21,1</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-26,-21,-21,-21</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-26,-5,-25,-5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-26,-15,-25,-15</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-26 0</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-439.5,52,-427</points>
<intersection>-439.5 2</intersection>
<intersection>-427 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-427,59,-427</points>
<connection>
<GID>780</GID>
<name>IN_6</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-439.5,52,-439.5</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,24,-29,25.5</points>
<intersection>24 3</intersection>
<intersection>25.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,25.5,-29,25.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,24,-28,24</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-435.5,53,-428</points>
<intersection>-435.5 2</intersection>
<intersection>-428 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-428,59,-428</points>
<connection>
<GID>780</GID>
<name>IN_5</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-435.5,53,-435.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,23,-29,23.5</points>
<intersection>23 3</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,23.5,-29,23.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,23,-28,23</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-431.5,54,-429</points>
<intersection>-431.5 2</intersection>
<intersection>-429 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-429,59,-429</points>
<connection>
<GID>780</GID>
<name>IN_4</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-431.5,54,-431.5</points>
<connection>
<GID>644</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,21.5,-29,22</points>
<intersection>21.5 2</intersection>
<intersection>22 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,21.5,-29,21.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,22,-28,22</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-430,55,-427.5</points>
<intersection>-430 1</intersection>
<intersection>-427.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-430,59,-430</points>
<connection>
<GID>780</GID>
<name>IN_3</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-427.5,55,-427.5</points>
<connection>
<GID>643</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,19.5,-29,21</points>
<intersection>19.5 2</intersection>
<intersection>21 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-30,19.5,-29,19.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,21,-28,21</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-431,56,-423.5</points>
<intersection>-431 1</intersection>
<intersection>-423.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-431,59,-431</points>
<connection>
<GID>780</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-423.5,56,-423.5</points>
<connection>
<GID>642</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,31,-32.5,32.5</points>
<intersection>31 1</intersection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,31,-28,31</points>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,32.5,-32.5,32.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-432,57,-419.5</points>
<intersection>-432 1</intersection>
<intersection>-419.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-432,59,-432</points>
<connection>
<GID>780</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-419.5,57,-419.5</points>
<connection>
<GID>641</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,30,-32.5,30.5</points>
<intersection>30 1</intersection>
<intersection>30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,30,-28,30</points>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,30.5,-32.5,30.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-433,58,-415.5</points>
<intersection>-433 1</intersection>
<intersection>-415.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-433,59,-433</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-415.5,58,-415.5</points>
<connection>
<GID>640</GID>
<name>OUT</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,28.5,-32.5,29</points>
<intersection>28.5 2</intersection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,29,-28,29</points>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,28.5,-32.5,28.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,26.5,-32.5,28</points>
<intersection>26.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,28,-28,28</points>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,26.5,-32.5,26.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39,-384,39,-384</points>
<connection>
<GID>784</GID>
<name>clock</name></connection>
<connection>
<GID>785</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-32,-78,-32</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39,-373,39,-373</points>
<connection>
<GID>784</GID>
<name>load</name></connection>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-34,-78,-34</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-392.5,28,-375</points>
<intersection>-392.5 2</intersection>
<intersection>-375 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-375,36,-375</points>
<connection>
<GID>784</GID>
<name>IN_7</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-392.5,28,-392.5</points>
<connection>
<GID>657</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-38,-78,-38</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-388.5,29,-376</points>
<intersection>-388.5 2</intersection>
<intersection>-376 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-376,36,-376</points>
<connection>
<GID>784</GID>
<name>IN_6</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-388.5,29,-388.5</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-36,-78,-36</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-384.5,30,-377</points>
<intersection>-384.5 2</intersection>
<intersection>-377 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-377,36,-377</points>
<connection>
<GID>784</GID>
<name>IN_5</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-384.5,30,-384.5</points>
<connection>
<GID>655</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-44,-78,-44</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-380.5,31,-378</points>
<intersection>-380.5 2</intersection>
<intersection>-378 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-378,36,-378</points>
<connection>
<GID>784</GID>
<name>IN_4</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-380.5,31,-380.5</points>
<connection>
<GID>654</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-42,-78,-42</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-379,32,-376.5</points>
<intersection>-379 1</intersection>
<intersection>-376.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-379,36,-379</points>
<connection>
<GID>784</GID>
<name>IN_3</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-376.5,32,-376.5</points>
<connection>
<GID>653</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-48,-78,-48</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-380,33,-372.5</points>
<intersection>-380 1</intersection>
<intersection>-372.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-380,36,-380</points>
<connection>
<GID>784</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-372.5,33,-372.5</points>
<connection>
<GID>652</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-46,-78,-46</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-381,34,-368.5</points>
<intersection>-381 1</intersection>
<intersection>-368.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-381,36,-381</points>
<connection>
<GID>784</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-368.5,34,-368.5</points>
<connection>
<GID>651</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,4,-33,12</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,12,-33,12</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-382,35,-364.5</points>
<intersection>-382 3</intersection>
<intersection>-364.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-364.5,35,-364.5</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-382,36,-382</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-460.5,43,-444.5</points>
<intersection>-460.5 2</intersection>
<intersection>-444.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,-460.5,43,-460.5</points>
<connection>
<GID>697</GID>
<name>OUT</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>43,-444.5,44,-444.5</points>
<connection>
<GID>647</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,4,-43,12</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,12,-43,12</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-43 0</intersection></hsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-456.5,42,-440.5</points>
<intersection>-456.5 2</intersection>
<intersection>-440.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-440.5,44,-440.5</points>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-456.5,42,-456.5</points>
<connection>
<GID>696</GID>
<name>OUT</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,4,-53,12</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,12,-53,12</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-53 0</intersection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-452.5,41,-436.5</points>
<intersection>-452.5 2</intersection>
<intersection>-436.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-436.5,44,-436.5</points>
<connection>
<GID>645</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-452.5,41,-452.5</points>
<connection>
<GID>695</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,4,-63,12</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,12,-63,12</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-448.5,40,-432.5</points>
<intersection>-448.5 2</intersection>
<intersection>-432.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-432.5,44,-432.5</points>
<connection>
<GID>644</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-448.5,40,-448.5</points>
<connection>
<GID>694</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-30,-63,-23</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-23,-63,-23</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-444.5,39,-428.5</points>
<intersection>-444.5 2</intersection>
<intersection>-428.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-428.5,44,-428.5</points>
<connection>
<GID>643</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-444.5,39,-444.5</points>
<connection>
<GID>693</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-30,-53,-23</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-23,-53,-23</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-53 0</intersection></hsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-440.5,38,-424.5</points>
<intersection>-440.5 2</intersection>
<intersection>-424.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-424.5,44,-424.5</points>
<connection>
<GID>642</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-440.5,38,-440.5</points>
<connection>
<GID>692</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-30,-43,-23</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-23,-43,-23</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-43 0</intersection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-436.5,37,-420.5</points>
<intersection>-436.5 2</intersection>
<intersection>-420.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-420.5,44,-420.5</points>
<connection>
<GID>641</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-436.5,37,-436.5</points>
<connection>
<GID>691</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-30,-33,-23</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-23,-33,-23</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-432.5,36,-416.5</points>
<intersection>-432.5 2</intersection>
<intersection>-416.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-416.5,44,-416.5</points>
<connection>
<GID>640</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-432.5,36,-432.5</points>
<connection>
<GID>689</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-27,69,-18.5</points>
<intersection>-27 2</intersection>
<intersection>-18.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,-27,69,-27</points>
<intersection>63 3</intersection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-27,63,-26</points>
<connection>
<GID>39</GID>
<name>A_greater_B</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>69,-18.5,71,-18.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-414.5,28,-398.5</points>
<intersection>-414.5 1</intersection>
<intersection>-398.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-414.5,44,-414.5</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-398.5,28,-398.5</points>
<connection>
<GID>666</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-45,70,-19.5</points>
<intersection>-45 2</intersection>
<intersection>-19.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,-45,70,-45</points>
<intersection>63 3</intersection>
<intersection>70 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-45,63,-44</points>
<connection>
<GID>49</GID>
<name>A_greater_B</name></connection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>70,-19.5,71,-19.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-418.5,29,-402.5</points>
<intersection>-418.5 1</intersection>
<intersection>-402.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-418.5,44,-418.5</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-402.5,29,-402.5</points>
<connection>
<GID>667</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-17.5,70,-9</points>
<intersection>-17.5 6</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,-9,70,-9</points>
<intersection>63 3</intersection>
<intersection>70 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-9,63,-8</points>
<connection>
<GID>54</GID>
<name>A_greater_B</name></connection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>70,-17.5,71,-17.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-422.5,30,-406.5</points>
<intersection>-422.5 1</intersection>
<intersection>-406.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-422.5,44,-422.5</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-406.5,30,-406.5</points>
<connection>
<GID>668</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-13.5,74,-11.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-426.5,31,-410.5</points>
<intersection>-426.5 1</intersection>
<intersection>-410.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-426.5,44,-426.5</points>
<connection>
<GID>643</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-410.5,31,-410.5</points>
<connection>
<GID>669</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-24.5,74,-22.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-430.5,32,-414.5</points>
<intersection>-430.5 1</intersection>
<intersection>-414.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-430.5,44,-430.5</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-414.5,32,-414.5</points>
<connection>
<GID>670</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-38,-2,-37,-2</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<connection>
<GID>77</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-434.5,33,-418.5</points>
<intersection>-434.5 1</intersection>
<intersection>-418.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-434.5,44,-434.5</points>
<connection>
<GID>645</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-418.5,33,-418.5</points>
<connection>
<GID>671</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-35,-2,-34,-2</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-438.5,34,-422.5</points>
<intersection>-438.5 1</intersection>
<intersection>-422.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-438.5,44,-438.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-422.5,34,-422.5</points>
<connection>
<GID>672</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-45,-2,-44,-2</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>75</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-442.5,35,-426.5</points>
<intersection>-442.5 1</intersection>
<intersection>-426.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-442.5,44,-442.5</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-426.5,35,-426.5</points>
<connection>
<GID>673</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-48,-2,-47,-2</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-420,-49,-393</points>
<intersection>-420 9</intersection>
<intersection>-407 12</intersection>
<intersection>-393 11</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-49,-420,-16,-420</points>
<intersection>-49 0</intersection>
<intersection>-16 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-16,-420,-16,-418</points>
<connection>
<GID>626</GID>
<name>clear</name></connection>
<intersection>-420 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-53,-393,-22,-393</points>
<connection>
<GID>609</GID>
<name>clear</name></connection>
<connection>
<GID>608</GID>
<name>clear</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-50,-407,-49,-407</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-55,-2,-54,-2</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-58,-2,-57,-2</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,-2,-64,-2</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-68,-2,-67,-2</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,-10,-66,-8</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66,-10,-64,-10</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-35,4,-35,4</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-45,4,-45,4</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-55,4,-55,4</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,4,-65,4</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61,-7.5,-61,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-7.5,-58,-7.5</points>
<intersection>-61 0</intersection>
<intersection>-58 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-58,-10,-58,-7.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-61,4,-59,4</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>-61 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-7.5,-51,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,-7.5,-48,-7.5</points>
<intersection>-51 0</intersection>
<intersection>-48 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-51,4,-49,4</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-51 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-48,-10,-48,-7.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41,-7.5,-41,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41,-7.5,-38,-7.5</points>
<intersection>-41 0</intersection>
<intersection>-38 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-38,-10,-38,-7.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-41,4,-39,4</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-41 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,4,-67,10</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,10,-35,10</points>
<intersection>-72 16</intersection>
<intersection>-67 0</intersection>
<intersection>-65 3</intersection>
<intersection>-57 5</intersection>
<intersection>-55 7</intersection>
<intersection>-47 9</intersection>
<intersection>-45 11</intersection>
<intersection>-37 13</intersection>
<intersection>-35 15</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-65,8,-65,10</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-57,4,-57,10</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-55,8,-55,10</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-47,4,-47,10</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-45,8,-45,10</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-37,4,-37,10</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-35,8,-35,10</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>10 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-72,-25,-72,10</points>
<intersection>-25 17</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-82,-25,-35,-25</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-72 16</intersection>
<intersection>-67 39</intersection>
<intersection>-65 22</intersection>
<intersection>-57 35</intersection>
<intersection>-55 26</intersection>
<intersection>-47 36</intersection>
<intersection>-45 30</intersection>
<intersection>-37 37</intersection>
<intersection>-35 34</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-65,-26,-65,-25</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-55,-26,-55,-25</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-45,-26,-45,-25</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-35,-26,-35,-25</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-57,-30,-57,-25</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>-47,-30,-47,-25</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>-37,-30,-37,-25</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>-67,-30,-67,-25</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-25 17</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-10,-56,-8</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-10,-54,-10</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-10,-46,-8</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,-10,-44,-10</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-10,-36,-8</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-10,-34,-10</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-38,-36,-37,-36</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-35,-36,-34,-36</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-45,-36,-44,-36</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-48,-36,-47,-36</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>95</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-55,-36,-54,-36</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>92</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-58,-36,-57,-36</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,-36,-64,-36</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-68,-36,-67,-36</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,-44,-66,-42</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66,-44,-64,-44</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-35,-30,-35,-30</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-45,-30,-45,-30</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-55,-30,-55,-30</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,-30,-65,-30</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61,-41.5,-61,-30</points>
<intersection>-41.5 1</intersection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-41.5,-58,-41.5</points>
<intersection>-61 0</intersection>
<intersection>-58 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-58,-44,-58,-41.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-61,-30,-59,-30</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>-61 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,-41.5,-51,-30</points>
<intersection>-41.5 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,-41.5,-48,-41.5</points>
<intersection>-51 0</intersection>
<intersection>-48 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-51,-30,-49,-30</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-51 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-48,-44,-48,-41.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41,-41.5,-41,-30</points>
<intersection>-41.5 1</intersection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41,-41.5,-38,-41.5</points>
<intersection>-41 0</intersection>
<intersection>-38 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-38,-44,-38,-41.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-41,-30,-39,-30</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>-41 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56,-44,-56,-42</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-44,-54,-44</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-56 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-44,-46,-42</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,-44,-44,-44</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-44,-36,-42</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-44,-34,-44</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-69,-30,-69,-30</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-69,4,-69,4</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-5,-21,-5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-11,43,-11</points>
<connection>
<GID>53</GID>
<name>IN_B_3</name></connection>
<intersection>3 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3,-11,3,-1</points>
<intersection>-11 1</intersection>
<intersection>-1 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>2,-1,4,-1</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>3 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-10,43,-10</points>
<connection>
<GID>53</GID>
<name>IN_B_2</name></connection>
<intersection>11 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>11,-10,11,-1</points>
<intersection>-10 1</intersection>
<intersection>-1 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>10,-1,12,-1</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>11 3</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-9,43,-9</points>
<connection>
<GID>53</GID>
<name>IN_B_1</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-9,19,-1</points>
<intersection>-9 1</intersection>
<intersection>-1 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>18,-1,20,-1</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-6,-1,-4,-1</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>119</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-17,4.5,-17</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>3.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>3.5,-25,3.5,-17</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,-17,12.5,-17</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>11.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>11.5,-25,11.5,-17</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-17,20.5,-17</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>19.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>19.5,-25,19.5,-17</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-6,-17,-4,-17</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-10,-27,3</points>
<intersection>-10 2</intersection>
<intersection>-3 3</intersection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,3,-21,3</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,-10,-27,-10</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27,-3,-21,-3</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-44,-27,-13</points>
<intersection>-44 2</intersection>
<intersection>-19 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,-13,-21,-13</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,-44,-27,-44</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-27,-19,-21,-19</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,0,-14,2</points>
<intersection>0 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,0,-12,0</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,2,-14,2</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-14,-14,-2</points>
<intersection>-14 2</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-2,-12,-2</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,-14,-14,-14</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-16,-13,-4</points>
<intersection>-16 5</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-15,-4,-13,-4</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>-13 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-13,-16,-12,-16</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-20,-14,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-18,-12,-18</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,-20,-14,-20</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-15,-21,-15</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-25,27.5,-17</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-17,27.5,-17</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-33,27.5,-29</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-33,26.5,-30</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>19.5,-30,19.5,-29</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-30,26.5,-30</points>
<intersection>19.5 1</intersection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-33,25.5,-31</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>11.5,-31,11.5,-29</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-31,25.5,-31</points>
<intersection>11.5 1</intersection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>3.5,-32,3.5,-29</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-32,24.5,-32</points>
<intersection>3.5 1</intersection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-33,24.5,-32</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>-32 2</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>34.5,-33,34.5,-33</points>
<connection>
<GID>1</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-41,39,-15</points>
<intersection>-41 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-15,43,-15</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-41,39,-41</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-42,40,-16</points>
<intersection>-42 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-16,43,-16</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-42,40,-42</points>
<intersection>30 3</intersection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-42,30,-41</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>-42 2</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-43,41,-17</points>
<intersection>-43 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-17,43,-17</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-43,41,-43</points>
<intersection>29 3</intersection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-43,29,-41</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-44,42,-18</points>
<intersection>-44 2</intersection>
<intersection>-18 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28,-44,42,-44</points>
<intersection>28 3</intersection>
<intersection>42 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-44,28,-41</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42,-18,43,-18</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-5,-52,-5,-4</points>
<intersection>-52 5</intersection>
<intersection>-24 45</intersection>
<intersection>-20 114</intersection>
<intersection>-8 44</intersection>
<intersection>-4 110</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-73,-52,-5,-52</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-71 33</intersection>
<intersection>-65 9</intersection>
<intersection>-55 8</intersection>
<intersection>-45 13</intersection>
<intersection>-35 36</intersection>
<intersection>-5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-55,-52,-55,-47</points>
<intersection>-52 5</intersection>
<intersection>-47 107</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-65,-52,-65,-47</points>
<intersection>-52 5</intersection>
<intersection>-47 106</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-45,-52,-45,-47</points>
<intersection>-52 5</intersection>
<intersection>-47 108</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-71,-18,-35,-18</points>
<intersection>-71 33</intersection>
<intersection>-65 24</intersection>
<intersection>-55 23</intersection>
<intersection>-45 28</intersection>
<intersection>-35 27</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-55,-18,-55,-13</points>
<intersection>-18 20</intersection>
<intersection>-13 103</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-65,-18,-65,-13</points>
<intersection>-18 20</intersection>
<intersection>-13 102</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>-35,-18,-35,-13</points>
<intersection>-18 20</intersection>
<intersection>-13 105</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-45,-18,-45,-13</points>
<intersection>-18 20</intersection>
<intersection>-13 104</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>-71,-52,-71,-18</points>
<intersection>-52 5</intersection>
<intersection>-18 20</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>-35,-52,-35,-47</points>
<intersection>-52 5</intersection>
<intersection>-47 109</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>-5,-8,20,-8</points>
<intersection>-5 3</intersection>
<intersection>4 81</intersection>
<intersection>12 85</intersection>
<intersection>20 87</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-5,-24,20.5,-24</points>
<intersection>-5 3</intersection>
<intersection>4.5 89</intersection>
<intersection>12.5 93</intersection>
<intersection>20.5 95</intersection></hsegment>
<vsegment>
<ID>81</ID>
<points>4,-8,4,-4</points>
<connection>
<GID>116</GID>
<name>clock</name></connection>
<intersection>-8 44</intersection></vsegment>
<vsegment>
<ID>85</ID>
<points>12,-8,12,-4</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<intersection>-8 44</intersection></vsegment>
<vsegment>
<ID>87</ID>
<points>20,-8,20,-4</points>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<intersection>-8 44</intersection></vsegment>
<vsegment>
<ID>89</ID>
<points>4.5,-24,4.5,-20</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>-24 45</intersection></vsegment>
<vsegment>
<ID>93</ID>
<points>12.5,-24,12.5,-20</points>
<connection>
<GID>122</GID>
<name>clock</name></connection>
<intersection>-24 45</intersection></vsegment>
<vsegment>
<ID>95</ID>
<points>20.5,-24,20.5,-20</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>-24 45</intersection></vsegment>
<hsegment>
<ID>102</ID>
<points>-65,-13,-64,-13</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>-65 24</intersection></hsegment>
<hsegment>
<ID>103</ID>
<points>-55,-13,-54,-13</points>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<intersection>-55 23</intersection></hsegment>
<hsegment>
<ID>104</ID>
<points>-45,-13,-44,-13</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>-45 28</intersection></hsegment>
<hsegment>
<ID>105</ID>
<points>-35,-13,-34,-13</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-35 27</intersection></hsegment>
<hsegment>
<ID>106</ID>
<points>-65,-47,-64,-47</points>
<connection>
<GID>88</GID>
<name>clock</name></connection>
<intersection>-65 9</intersection></hsegment>
<hsegment>
<ID>107</ID>
<points>-55,-47,-54,-47</points>
<connection>
<GID>94</GID>
<name>clock</name></connection>
<intersection>-55 8</intersection></hsegment>
<hsegment>
<ID>108</ID>
<points>-45,-47,-44,-47</points>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<intersection>-45 13</intersection></hsegment>
<hsegment>
<ID>109</ID>
<points>-35,-47,-34,-47</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<intersection>-35 36</intersection></hsegment>
<hsegment>
<ID>110</ID>
<points>-5,-4,-4,-4</points>
<connection>
<GID>115</GID>
<name>clock</name></connection>
<intersection>-5 3</intersection></hsegment>
<hsegment>
<ID>114</ID>
<points>-5,-20,-4,-20</points>
<connection>
<GID>120</GID>
<name>clock</name></connection>
<intersection>-5 3</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,5,60,6.5</points>
<intersection>5 3</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,6.5,60,6.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,5,61,5</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,4.5,61,4.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>61 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>61,4,61,4.5</points>
<connection>
<GID>54</GID>
<name>IN_B_1</name></connection>
<intersection>4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,2.5,60,3</points>
<intersection>2.5 2</intersection>
<intersection>3 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,2.5,60,2.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,3,61,3</points>
<connection>
<GID>54</GID>
<name>IN_B_2</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,0.5,60,2</points>
<intersection>0.5 2</intersection>
<intersection>2 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,0.5,60,0.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,2,61,2</points>
<connection>
<GID>54</GID>
<name>IN_B_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-13,60,-11.5</points>
<intersection>-13 3</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-11.5,60,-11.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-13,61,-13</points>
<connection>
<GID>39</GID>
<name>IN_B_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-14,60,-13.5</points>
<intersection>-14 3</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-13.5,60,-13.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-14,61,-14</points>
<connection>
<GID>39</GID>
<name>IN_B_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-15.5,60,-15</points>
<intersection>-15.5 2</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-15.5,60,-15.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-15,61,-15</points>
<connection>
<GID>39</GID>
<name>IN_B_2</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-17.5,60,-16</points>
<intersection>-17.5 2</intersection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-17.5,60,-17.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-16,61,-16</points>
<connection>
<GID>39</GID>
<name>IN_B_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-31,60,-29.5</points>
<intersection>-31 3</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-29.5,60,-29.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-31,61,-31</points>
<connection>
<GID>49</GID>
<name>IN_B_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-32,60,-31.5</points>
<intersection>-32 3</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-31.5,60,-31.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-32,61,-32</points>
<connection>
<GID>49</GID>
<name>IN_B_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-33.5,60,-33</points>
<intersection>-33.5 2</intersection>
<intersection>-33 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-33.5,60,-33.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-33,61,-33</points>
<connection>
<GID>49</GID>
<name>IN_B_2</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-35.5,60,-34</points>
<intersection>-35.5 2</intersection>
<intersection>-34 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-35.5,60,-35.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-34,61,-34</points>
<connection>
<GID>49</GID>
<name>IN_B_3</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-2,61,-2</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>52 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52,-38,52,-2</points>
<intersection>-38 7</intersection>
<intersection>-20 5</intersection>
<intersection>-11.5 8</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>52,-20,61,-20</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>52 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>52,-38,61,-38</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>52 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>51,-11.5,52,-11.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>52 3</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-39,53,-3</points>
<intersection>-39 5</intersection>
<intersection>-21 3</intersection>
<intersection>-12.5 2</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-3,61,-3</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-12.5,53,-12.5</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,-21,61,-21</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>53,-39,61,-39</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-40,54,-4</points>
<intersection>-40 5</intersection>
<intersection>-22 3</intersection>
<intersection>-13.5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-4,61,-4</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-13.5,54,-13.5</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54,-22,61,-22</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54,-40,61,-40</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-41,55,-5</points>
<intersection>-41 5</intersection>
<intersection>-23 3</intersection>
<intersection>-14.5 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-5,61,-5</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-14.5,55,-14.5</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>55,-23,61,-23</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>55,-41,61,-41</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-8,43,-8</points>
<connection>
<GID>53</GID>
<name>IN_B_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-8,27,-1</points>
<intersection>-8 1</intersection>
<intersection>-1 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26,-1,27,-1</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>27 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-99.5,-7.5,-95.5</points>
<intersection>-99.5 4</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-95.5,-7.5,-95.5</points>
<intersection>-15.5 3</intersection>
<intersection>-7.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15.5,-95.5,-15.5,-93.5</points>
<intersection>-95.5 2</intersection>
<intersection>-93.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-8.5,-99.5,-6.5,-99.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-15.5,-93.5,-14.5,-93.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-96.5,-8.5,-96.5</points>
<intersection>-14.5 3</intersection>
<intersection>-8.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-98.5,-14.5,-96.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-8.5,-96.5,-8.5,-92.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>-96.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-102,-51.5,-100.5</points>
<intersection>-102 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-100.5,-50.5,-100.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-102,-51.5,-102</points>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-103,-51.5,-102.5</points>
<intersection>-103 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-102.5,-50.5,-102.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-103,-51.5,-103</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-104.5,-51.5,-104</points>
<intersection>-104.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-104.5,-50.5,-104.5</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-104,-51.5,-104</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-106.5,-51.5,-105</points>
<intersection>-106.5 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-106.5,-50.5,-106.5</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-105,-51.5,-105</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-99,-26.5,-84</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-99 6</intersection>
<intersection>-95 3</intersection>
<intersection>-85.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-26.5,-95,-22.5,-95</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-26.5,-99,-22.5,-99</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-26.5,-85.5,-24.5,-85.5</points>
<intersection>-26.5 0</intersection>
<intersection>-24.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-24.5,-86,-24.5,-85.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-85.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-110,-57.5,-108</points>
<connection>
<GID>129</GID>
<name>clock</name></connection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-110,-57.5,-110</points>
<connection>
<GID>132</GID>
<name>CLK</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-104,-62.5,-100</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>-100 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,-100,-62.5,-100</points>
<intersection>-68.5 3</intersection>
<intersection>-62.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68.5,-100,-68.5,-98</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>-100 2</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-101,-61.5,-101</points>
<intersection>-69.5 3</intersection>
<intersection>-61.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-69.5,-103,-69.5,-101</points>
<intersection>-103 17</intersection>
<intersection>-101 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-61.5,-101,-61.5,-97</points>
<intersection>-101 1</intersection>
<intersection>-97 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-62.5,-97,-56.5,-97</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>-61.5 4</intersection>
<intersection>-56.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-56.5,-99,-56.5,-97</points>
<connection>
<GID>129</GID>
<name>count_enable</name></connection>
<intersection>-97 15</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-69.5,-103,-68.5,-103</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-69.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-104,-34.5,-100</points>
<intersection>-104 2</intersection>
<intersection>-100 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-104,-34.5,-104</points>
<intersection>-40.5 3</intersection>
<intersection>-34.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40.5,-106,-40.5,-104</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-34.5,-100,-28.5,-100</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>-34.5 0</intersection>
<intersection>-32.5 12</intersection>
<intersection>-28.5 8</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-28.5,-97,-22.5,-97</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-28.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-28.5,-110,-28.5,-97</points>
<intersection>-110 9</intersection>
<intersection>-100 4</intersection>
<intersection>-97 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-28.5,-110,-22.5,-110</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-28.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-32.5,-117,-32.5,-100</points>
<intersection>-117 13</intersection>
<intersection>-100 4</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-75.5,-117,-32.5,-117</points>
<intersection>-75.5 14</intersection>
<intersection>-54.5 17</intersection>
<intersection>-32.5 12</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-75.5,-117,-75.5,-97</points>
<intersection>-117 13</intersection>
<intersection>-97 18</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>-54.5,-117,-54.5,-116</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>-117 13</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-75.5,-97,-74.5,-97</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>-75.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-108,-42.5,-103.5</points>
<intersection>-108 1</intersection>
<intersection>-103.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42.5,-108,-40.5,-108</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-103.5,-42.5,-103.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-107,-33.5,-103</points>
<intersection>-107 4</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-41.5,-103,-33.5,-103</points>
<intersection>-41.5 3</intersection>
<intersection>-33.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-41.5,-103,-41.5,-101</points>
<intersection>-103 2</intersection>
<intersection>-101 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-34.5,-107,-33.5,-107</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-41.5,-101,-40.5,-101</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>-41.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-70.5,-105,-68.5,-105</points>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,-96,-68.5,-96</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-110,-55.5,-108</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-94,-16.5,-91.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-91.5,-14.5,-91.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-100.5,-16.5,-98</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,-100.5,-14.5,-100.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-112.5,-7.5,-108.5</points>
<intersection>-112.5 4</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-108.5,-7.5,-108.5</points>
<intersection>-15.5 3</intersection>
<intersection>-7.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15.5,-108.5,-15.5,-106.5</points>
<intersection>-108.5 2</intersection>
<intersection>-106.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-8.5,-112.5,-6.5,-112.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-15.5,-106.5,-14.5,-106.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>-15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-109.5,-8.5,-109.5</points>
<intersection>-14.5 3</intersection>
<intersection>-8.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-111.5,-14.5,-109.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>-109.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-8.5,-109.5,-8.5,-105.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>-109.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-107,-16.5,-104.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16.5,-104.5,-14.5,-104.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16.5,-113.5,-16.5,-111</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,-113.5,-14.5,-113.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>-16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-112,-24.5,-90</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-108,-22.5,-108</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-24.5,-112,-22.5,-112</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-78.5,-93,-22.5,-93</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-76.5 8</intersection>
<intersection>-75.5 20</intersection>
<intersection>-42.5 5</intersection>
<intersection>-30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30.5,-106,-30.5,-93</points>
<intersection>-106 4</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-30.5,-106,-22.5,-106</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-30.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-42.5,-99,-42.5,-93</points>
<intersection>-99 32</intersection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-76.5,-118,-76.5,-93</points>
<intersection>-118 21</intersection>
<intersection>-105 18</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-76.5,-105,-74.5,-105</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-76.5 8</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-75.5,-95,-75.5,-93</points>
<intersection>-95 33</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-76.5,-118,-56.5,-118</points>
<intersection>-76.5 8</intersection>
<intersection>-56.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-56.5,-118,-56.5,-116</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-118 21</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>-42.5,-99,-40.5,-99</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-42.5 5</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>-75.5,-95,-74.5,-95</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-75.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-181.5,49.5,-181.5</points>
<connection>
<GID>159</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-189.5,49.5,-189.5</points>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<connection>
<GID>162</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-197.5,49.5,-197.5</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<connection>
<GID>164</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-205.5,49.5,-205.5</points>
<connection>
<GID>165</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>49.5,-213.5,49.5,-213.5</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-221.5,49.5,-221.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<connection>
<GID>170</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-229.5,49.5,-229.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<connection>
<GID>172</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-237.5,49.5,-237.5</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-232.5,38.5,-172.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>-232.5 13</intersection>
<intersection>-216.5 10</intersection>
<intersection>-200.5 5</intersection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-184.5,43.5,-184.5</points>
<connection>
<GID>160</GID>
<name>IN_3</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-200.5,43.5,-200.5</points>
<connection>
<GID>164</GID>
<name>IN_3</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>38.5,-216.5,43.5,-216.5</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>38.5,-232.5,43.5,-232.5</points>
<connection>
<GID>172</GID>
<name>IN_3</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-222.5,35,-172.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-222.5 16</intersection>
<intersection>-214.5 11</intersection>
<intersection>-190.5 3</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-182.5,43.5,-182.5</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-190.5,43.5,-190.5</points>
<connection>
<GID>162</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>35,-214.5,43.5,-214.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>35,-222.5,43.5,-222.5</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-204.5,31.5,-172.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>-204.5 7</intersection>
<intersection>-196.5 5</intersection>
<intersection>-188.5 3</intersection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-180.5,43.5,-180.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31.5,-188.5,43.5,-188.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31.5,-196.5,43.5,-196.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31.5,-204.5,43.5,-204.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-178.5,43.5,-178.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>15.5 29</intersection>
<intersection>23 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>23,-234.5,23,-178.5</points>
<intersection>-234.5 15</intersection>
<intersection>-226.5 17</intersection>
<intersection>-218.5 18</intersection>
<intersection>-210.5 19</intersection>
<intersection>-202.5 20</intersection>
<intersection>-194.5 21</intersection>
<intersection>-186.5 16</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>23,-234.5,43.5,-234.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>23,-186.5,43.5,-186.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>23,-226.5,43.5,-226.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>23,-218.5,43.5,-218.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>23,-210.5,43.5,-210.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>23,-202.5,43.5,-202.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>23,-194.5,43.5,-194.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>23 13</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>15.5,-203,15.5,-178.5</points>
<intersection>-203 30</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>13,-203,15.5,-203</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>15.5 29</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>20</ID>
<points>-84,-168.5,234.5,-168.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>37 21</intersection>
<intersection>40.5 32</intersection>
<intersection>234.5 31</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>37,-224.5,37,-168.5</points>
<intersection>-224.5 27</intersection>
<intersection>-208.5 26</intersection>
<intersection>-192.5 25</intersection>
<intersection>-168.5 20</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>37,-192.5,43.5,-192.5</points>
<connection>
<GID>162</GID>
<name>IN_3</name></connection>
<intersection>37 21</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>37,-208.5,43.5,-208.5</points>
<connection>
<GID>166</GID>
<name>IN_3</name></connection>
<intersection>37 21</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>37,-224.5,43.5,-224.5</points>
<connection>
<GID>170</GID>
<name>IN_3</name></connection>
<intersection>37 21</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>234.5,-257,234.5,-168.5</points>
<connection>
<GID>256</GID>
<name>SEL_0</name></connection>
<intersection>-168.5 20</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>40.5,-240.5,40.5,-168.5</points>
<intersection>-240.5 33</intersection>
<intersection>-168.5 20</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>40.5,-240.5,43.5,-240.5</points>
<connection>
<GID>174</GID>
<name>IN_3</name></connection>
<intersection>40.5 32</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>23</ID>
<points>-84,-166.5,233.5,-166.5</points>
<connection>
<GID>395</GID>
<name>OUT_0</name></connection>
<intersection>33.5 24</intersection>
<intersection>35 36</intersection>
<intersection>233.5 37</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>33.5,-238.5,33.5,-166.5</points>
<intersection>-238.5 39</intersection>
<intersection>-230.5 32</intersection>
<intersection>-206.5 30</intersection>
<intersection>-198.5 28</intersection>
<intersection>-166.5 23</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>33.5,-198.5,43.5,-198.5</points>
<connection>
<GID>164</GID>
<name>IN_2</name></connection>
<intersection>33.5 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>33.5,-206.5,43.5,-206.5</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>33.5 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>33.5,-230.5,43.5,-230.5</points>
<connection>
<GID>172</GID>
<name>IN_2</name></connection>
<intersection>33.5 24</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>35,-168.5,35,-166.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>-166.5 23</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>233.5,-257,233.5,-166.5</points>
<connection>
<GID>256</GID>
<name>SEL_1</name></connection>
<intersection>-166.5 23</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>33.5,-238.5,43.5,-238.5</points>
<connection>
<GID>174</GID>
<name>IN_2</name></connection>
<intersection>33.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>22</ID>
<points>-84,-164.5,232.5,-164.5</points>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection>
<intersection>30 23</intersection>
<intersection>31.5 36</intersection>
<intersection>232.5 37</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>30,-236.5,30,-164.5</points>
<intersection>-236.5 39</intersection>
<intersection>-228.5 31</intersection>
<intersection>-220.5 29</intersection>
<intersection>-212.5 27</intersection>
<intersection>-164.5 22</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>30,-212.5,43.5,-212.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>30 23</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>30,-220.5,43.5,-220.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>30 23</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>30,-228.5,43.5,-228.5</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>30 23</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>31.5,-168.5,31.5,-164.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-164.5 22</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>232.5,-257,232.5,-164.5</points>
<connection>
<GID>256</GID>
<name>SEL_2</name></connection>
<intersection>-164.5 22</intersection></vsegment>
<hsegment>
<ID>39</ID>
<points>30,-236.5,43.5,-236.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>30 23</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-51,-195,-50,-195</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<connection>
<GID>180</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-48,-195,-47,-195</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>19</ID>
<points>18,-219,18,-174</points>
<intersection>-219 79</intersection>
<intersection>-174 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>18,-174,143.5,-174</points>
<intersection>18 19</intersection>
<intersection>143.5 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>143.5,-274,143.5,-174</points>
<intersection>-274 47</intersection>
<intersection>-214 69</intersection>
<intersection>-174 24</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>143.5,-274,214.5,-274</points>
<intersection>143.5 36</intersection>
<intersection>160 77</intersection>
<intersection>169 59</intersection>
<intersection>178 60</intersection>
<intersection>187.5 61</intersection>
<intersection>196.5 63</intersection>
<intersection>205.5 64</intersection>
<intersection>214.5 65</intersection></hsegment>
<vsegment>
<ID>59</ID>
<points>169,-274.5,169,-274</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<vsegment>
<ID>60</ID>
<points>178,-274.5,178,-274</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>187.5,-274.5,187.5,-274</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>196.5,-274.5,196.5,-274</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>205.5,-274.5,205.5,-274</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<vsegment>
<ID>65</ID>
<points>214.5,-274.5,214.5,-274</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<hsegment>
<ID>69</ID>
<points>143.5,-214,213,-214</points>
<intersection>143.5 36</intersection>
<intersection>158.5 76</intersection>
<intersection>167.5 75</intersection>
<intersection>176.5 74</intersection>
<intersection>186 73</intersection>
<intersection>195 72</intersection>
<intersection>204 71</intersection>
<intersection>213 70</intersection></hsegment>
<vsegment>
<ID>70</ID>
<points>213,-215,213,-214</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>71</ID>
<points>204,-215,204,-214</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>72</ID>
<points>195,-215,195,-214</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>186,-215,186,-214</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>176.5,-215,176.5,-214</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>167.5,-215,167.5,-214</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>158.5,-215,158.5,-214</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-214 69</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>160,-274.5,160,-274</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-274 47</intersection></vsegment>
<hsegment>
<ID>79</ID>
<points>-29,-219,18,-219</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>18 19</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-200.5,-53.5,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53.5,-200.5,-50.5,-200.5</points>
<intersection>-53.5 0</intersection>
<intersection>-50.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-189,-52,-189</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-50.5,-203,-50.5,-200.5</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-42,-195,-41,-195</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<connection>
<GID>189</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-39,-195,-38,-195</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-200.5,-44.5,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-200.5,-41.5,-200.5</points>
<intersection>-44.5 0</intersection>
<intersection>-41.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44.5,-189,-43,-189</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-41.5,-203,-41.5,-200.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-33,-195,-32,-195</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>193</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-30,-195,-29,-195</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<connection>
<GID>194</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-200.5,-35.5,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-200.5,-32.5,-200.5</points>
<intersection>-35.5 0</intersection>
<intersection>-32.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-35.5,-189,-34,-189</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-32.5,-203,-32.5,-200.5</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-23.5,-195,-22.5,-195</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<connection>
<GID>197</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-20.5,-195,-19.5,-195</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>198</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-200.5,-26,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-200.5,-23,-200.5</points>
<intersection>-26 0</intersection>
<intersection>-23 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,-189,-24.5,-189</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>-26 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-23,-203,-23,-200.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-14.5,-195,-13.5,-195</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>201</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-11.5,-195,-10.5,-195</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,-200.5,-17,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,-200.5,-14,-200.5</points>
<intersection>-17 0</intersection>
<intersection>-14 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17,-189,-15.5,-189</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>-17 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14,-203,-14,-200.5</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-5.5,-195,-4.5,-195</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<connection>
<GID>205</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2.5,-195,-1.5,-195</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-200.5,-8,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-200.5,-5,-200.5</points>
<intersection>-8 0</intersection>
<intersection>-5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-189,-6.5,-189</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>-8 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-5,-203,-5,-200.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>3.5,-195,4.5,-195</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>209</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>6.5,-195,7.5,-195</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-200.5,1,-189</points>
<intersection>-200.5 1</intersection>
<intersection>-189 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-200.5,4,-200.5</points>
<intersection>1 0</intersection>
<intersection>4 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-189,2.5,-189</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>1 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4,-203,4,-200.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,-203,-59,-185.5</points>
<intersection>-203 4</intersection>
<intersection>-185.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-62.5,-185.5,-59,-185.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>-59 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-59,-203,-56.5,-203</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,-189,-48,-184.5</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-184.5,-48,-184.5</points>
<connection>
<GID>213</GID>
<name>OUT_1</name></connection>
<intersection>-48 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-203,-49,-201</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-203,-47.5,-203</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-203,-31,-201</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31,-203,-29,-203</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-203,-40,-201</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-203,-38.5,-203</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-40 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-203,-21.5,-201</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-203,-20,-203</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-203,-12.5,-201</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-203,-11,-203</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-203,-3.5,-201</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-203,-2,-203</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-203,5.5,-201</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>-203 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-203,7,-203</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-189,6.5,-178.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-178.5,6.5,-178.5</points>
<connection>
<GID>213</GID>
<name>OUT_7</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-189,-2.5,-179.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>-179.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-179.5,-2.5,-179.5</points>
<connection>
<GID>213</GID>
<name>OUT_6</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-189,-11.5,-180.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>-180.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-180.5,-11.5,-180.5</points>
<connection>
<GID>213</GID>
<name>OUT_5</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-189,-20.5,-181.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>-181.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-181.5,-20.5,-181.5</points>
<connection>
<GID>213</GID>
<name>OUT_4</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-189,-30,-182.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-182.5,-30,-182.5</points>
<connection>
<GID>213</GID>
<name>OUT_3</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-189,-39,-183.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>-183.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,-183.5,-39,-183.5</points>
<connection>
<GID>213</GID>
<name>OUT_2</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>58</ID>
<points>-39,-250,125.5,-250</points>
<intersection>-39 1038</intersection>
<intersection>125.5 148</intersection></hsegment>
<hsegment>
<ID>110</ID>
<points>125.5,-254,211.5,-254</points>
<intersection>125.5 148</intersection>
<intersection>148 1011</intersection>
<intersection>157 1012</intersection>
<intersection>166 1013</intersection>
<intersection>175.5 1014</intersection>
<intersection>184.5 1015</intersection>
<intersection>193.5 1016</intersection>
<intersection>202.5 1017</intersection>
<intersection>211.5 1018</intersection></hsegment>
<vsegment>
<ID>148</ID>
<points>125.5,-309,125.5,-250</points>
<intersection>-309 150</intersection>
<intersection>-254 110</intersection>
<intersection>-250 58</intersection></vsegment>
<hsegment>
<ID>150</ID>
<points>125.5,-309,213,-309</points>
<intersection>125.5 148</intersection>
<intersection>149.5 1019</intersection>
<intersection>158.5 1020</intersection>
<intersection>167.5 1021</intersection>
<intersection>177 1022</intersection>
<intersection>186 1023</intersection>
<intersection>195 1024</intersection>
<intersection>204 1025</intersection>
<intersection>213 180</intersection></hsegment>
<vsegment>
<ID>180</ID>
<points>213,-330,213,-291.5</points>
<connection>
<GID>291</GID>
<name>clock</name></connection>
<intersection>-330 235</intersection>
<intersection>-309 150</intersection></vsegment>
<hsegment>
<ID>235</ID>
<points>213,-330,361.5,-330</points>
<intersection>213 180</intersection>
<intersection>361.5 1040</intersection></hsegment>
<vsegment>
<ID>1011</ID>
<points>148,-254,148,-232</points>
<connection>
<GID>294</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1012</ID>
<points>157,-254,157,-232</points>
<connection>
<GID>302</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1013</ID>
<points>166,-254,166,-232</points>
<connection>
<GID>307</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1014</ID>
<points>175.5,-254,175.5,-232</points>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1015</ID>
<points>184.5,-254,184.5,-232</points>
<connection>
<GID>315</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1016</ID>
<points>193.5,-254,193.5,-232</points>
<connection>
<GID>319</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1017</ID>
<points>202.5,-254,202.5,-232</points>
<connection>
<GID>323</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1018</ID>
<points>211.5,-254,211.5,-232</points>
<connection>
<GID>327</GID>
<name>clock</name></connection>
<intersection>-254 110</intersection></vsegment>
<vsegment>
<ID>1019</ID>
<points>149.5,-309,149.5,-291.5</points>
<connection>
<GID>261</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1020</ID>
<points>158.5,-309,158.5,-291.5</points>
<connection>
<GID>267</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1021</ID>
<points>167.5,-309,167.5,-291.5</points>
<connection>
<GID>271</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1022</ID>
<points>177,-309,177,-291.5</points>
<connection>
<GID>275</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1023</ID>
<points>186,-309,186,-291.5</points>
<connection>
<GID>279</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1024</ID>
<points>195,-309,195,-291.5</points>
<connection>
<GID>283</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1025</ID>
<points>204,-309,204,-291.5</points>
<connection>
<GID>287</GID>
<name>clock</name></connection>
<intersection>-309 150</intersection></vsegment>
<vsegment>
<ID>1038</ID>
<points>-39,-250,-39,-236</points>
<intersection>-250 58</intersection>
<intersection>-236 1039</intersection></vsegment>
<hsegment>
<ID>1039</ID>
<points>-54,-236,-39,-236</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>-39 1038</intersection></hsegment>
<vsegment>
<ID>1040</ID>
<points>361.5,-330,361.5,-303.5</points>
<intersection>-330 235</intersection>
<intersection>-303.5 1041</intersection></vsegment>
<hsegment>
<ID>1041</ID>
<points>361.5,-303.5,365.5,-303.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>361.5 1040</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-82.5,-227.5,-80,-227.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-82.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-82.5,-229,-82.5,-227.5</points>
<intersection>-229 12</intersection>
<intersection>-227.5 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-88.5,-229,-82.5,-229</points>
<connection>
<GID>214</GID>
<name>CLK</name></connection>
<intersection>-82.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,-223.5,-86.5,-223.5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<connection>
<GID>219</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,-225.5,-80,-224.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-224.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-80.5,-224.5,-80,-224.5</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>-80 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,-225.5,-86.5,-225.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-94 14</intersection>
<intersection>-88 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88,-231,-88,-225.5</points>
<intersection>-231 16</intersection>
<intersection>-225.5 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>-94,-225.5,-94,-220</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-88,-231,-81.5,-231</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-88 9</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,-231,-70.5,-226.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,-231,-70.5,-231</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-74.5,-219.5,-71.5,-219.5</points>
<connection>
<GID>216</GID>
<name>clock</name></connection>
<intersection>-71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71.5,-220.5,-71.5,-219.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>-219.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-83.5,-218.5,-83.5,-218.5</points>
<connection>
<GID>216</GID>
<name>count_enable</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90.5,-223.5,-90.5,-207.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-207.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-90.5,-207.5,-74.5,-207.5</points>
<intersection>-90.5 0</intersection>
<intersection>-79 3</intersection>
<intersection>-74.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-74.5,-217.5,-74.5,-207.5</points>
<connection>
<GID>216</GID>
<name>clear</name></connection>
<intersection>-207.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-79,-208,-79,-207.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>-207.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,-214.5,-80.5,-214</points>
<connection>
<GID>216</GID>
<name>OUT_3</name></connection>
<intersection>-214 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-80.5,-214,-80,-214</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-237,84.5,-237</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>70 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>70,-237,70,-181.5</points>
<intersection>-237 1</intersection>
<intersection>-181.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>51.5,-181.5,70,-181.5</points>
<connection>
<GID>159</GID>
<name>N_in1</name></connection>
<intersection>70 2</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-231,84.5,-209.5</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>-209.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-209.5,107.5,-209.5</points>
<intersection>84.5 0</intersection>
<intersection>107.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>107.5,-211,107.5,-209.5</points>
<intersection>-211 3</intersection>
<intersection>-209.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-211,109.5,-211</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>107.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-222.5,84.5,-200.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-200.5,106.5,-200.5</points>
<intersection>84.5 0</intersection>
<intersection>106.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>106.5,-210,106.5,-200.5</points>
<intersection>-210 5</intersection>
<intersection>-200.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>106.5,-210,109.5,-210</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>106.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-214,84.5,-192</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-192 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-192,105.5,-192</points>
<intersection>84.5 0</intersection>
<intersection>105.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>105.5,-209,105.5,-192</points>
<intersection>-209 8</intersection>
<intersection>-192 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>105.5,-209,109.5,-209</points>
<connection>
<GID>220</GID>
<name>IN_2</name></connection>
<intersection>105.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-206,84.5,-184</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-184 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-184,104.5,-184</points>
<intersection>84.5 0</intersection>
<intersection>104.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>104.5,-208,104.5,-184</points>
<intersection>-208 5</intersection>
<intersection>-184 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>104.5,-208,109.5,-208</points>
<connection>
<GID>220</GID>
<name>IN_3</name></connection>
<intersection>104.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-207,105.5,-197.5</points>
<intersection>-207 5</intersection>
<intersection>-197.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>105.5,-207,109.5,-207</points>
<connection>
<GID>220</GID>
<name>IN_4</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-197.5,105.5,-197.5</points>
<intersection>84.5 8</intersection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>84.5,-198.5,84.5,-197</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>-197.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-191,84.5,-169</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-169 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-169,106.5,-169</points>
<intersection>84.5 0</intersection>
<intersection>106.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>106.5,-206,106.5,-169</points>
<intersection>-206 5</intersection>
<intersection>-169 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>106.5,-206,109.5,-206</points>
<connection>
<GID>220</GID>
<name>IN_5</name></connection>
<intersection>106.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-183.5,84.5,-161.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>-161.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-161.5,107.5,-161.5</points>
<intersection>84.5 0</intersection>
<intersection>107.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>107.5,-205,107.5,-161.5</points>
<intersection>-205 5</intersection>
<intersection>-161.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>107.5,-205,109.5,-205</points>
<connection>
<GID>220</GID>
<name>IN_6</name></connection>
<intersection>107.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-176,84.5,-175.5</points>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection>
<intersection>-175.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-175.5,109.5,-175.5</points>
<intersection>84.5 0</intersection>
<intersection>109.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>109.5,-204,109.5,-175.5</points>
<connection>
<GID>220</GID>
<name>IN_7</name></connection>
<intersection>-175.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-202,112.5,-202</points>
<connection>
<GID>220</GID>
<name>load</name></connection>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-321,67,-189.5</points>
<intersection>-321 3</intersection>
<intersection>-189.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-189.5,67,-189.5</points>
<connection>
<GID>161</GID>
<name>N_in1</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67,-321,86.5,-321</points>
<intersection>67 0</intersection>
<intersection>86.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>86.5,-321,86.5,-320</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-321 3</intersection></vsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-314,86.5,-292.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>-292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-292.5,109.5,-292.5</points>
<intersection>86.5 0</intersection>
<intersection>109.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>109.5,-294,109.5,-292.5</points>
<intersection>-294 3</intersection>
<intersection>-292.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>109.5,-294,111.5,-294</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>109.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-305.5,86.5,-284</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-284 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-284,108.5,-284</points>
<intersection>86.5 0</intersection>
<intersection>108.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>108.5,-293,108.5,-284</points>
<intersection>-293 5</intersection>
<intersection>-284 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>108.5,-293,111.5,-293</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>108.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-297,86.5,-275</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-275 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>86.5,-275,107.5,-275</points>
<intersection>86.5 0</intersection>
<intersection>107.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>107.5,-292,107.5,-275</points>
<intersection>-292 8</intersection>
<intersection>-275 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>107.5,-292,111.5,-292</points>
<connection>
<GID>230</GID>
<name>IN_2</name></connection>
<intersection>107.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-289,86.5,-267</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-267 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-267,106.5,-267</points>
<intersection>86.5 0</intersection>
<intersection>106.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>106.5,-291,106.5,-267</points>
<intersection>-291 5</intersection>
<intersection>-267 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>106.5,-291,111.5,-291</points>
<connection>
<GID>230</GID>
<name>IN_3</name></connection>
<intersection>106.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-290,107.5,-281</points>
<intersection>-290 5</intersection>
<intersection>-281 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>107.5,-290,111.5,-290</points>
<connection>
<GID>230</GID>
<name>IN_4</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>86.5,-281,107.5,-281</points>
<intersection>86.5 8</intersection>
<intersection>107.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>86.5,-281.5,86.5,-280</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-281 6</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-274,86.5,-252</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>-252 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-252,108.5,-252</points>
<intersection>86.5 0</intersection>
<intersection>108.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>108.5,-289,108.5,-252</points>
<intersection>-289 5</intersection>
<intersection>-252 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>108.5,-289,111.5,-289</points>
<connection>
<GID>230</GID>
<name>IN_5</name></connection>
<intersection>108.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-266.5,86.5,-244.5</points>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>86.5,-244.5,109.5,-244.5</points>
<intersection>86.5 0</intersection>
<intersection>109.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>109.5,-288,109.5,-244.5</points>
<intersection>-288 5</intersection>
<intersection>-244.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>109.5,-288,111.5,-288</points>
<connection>
<GID>230</GID>
<name>IN_6</name></connection>
<intersection>109.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-259,86.5,-256.5</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-256.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-256.5,111.5,-256.5</points>
<intersection>86.5 0</intersection>
<intersection>111.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>111.5,-287,111.5,-256.5</points>
<connection>
<GID>230</GID>
<name>IN_7</name></connection>
<intersection>-256.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-78.5,-206.5,-63,-206.5</points>
<intersection>-78.5 7</intersection>
<intersection>-63 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-63,-223.5,-63,-206.5</points>
<intersection>-223.5 5</intersection>
<intersection>-206.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-63,-223.5,-50.5,-223.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>-63 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-78.5,-206.5,-78.5,-204</points>
<intersection>-206.5 1</intersection>
<intersection>-204 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-80.5,-204,-77.5,-204</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>-78.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-285,114.5,-285</points>
<connection>
<GID>230</GID>
<name>load</name></connection>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,-178.5,-76.5,-176.5</points>
<intersection>-178.5 1</intersection>
<intersection>-176.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,-178.5,-70.5,-178.5</points>
<connection>
<GID>213</GID>
<name>IN_7</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-176.5,-76.5,-176.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-179.5,-77.5,-178.5</points>
<intersection>-179.5 2</intersection>
<intersection>-178.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83.5,-178.5,-77.5,-178.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77.5,-179.5,-70.5,-179.5</points>
<connection>
<GID>213</GID>
<name>IN_6</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-180.5,-70.5,-180.5</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,-182.5,-78,-181.5</points>
<intersection>-182.5 1</intersection>
<intersection>-181.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83.5,-182.5,-78,-182.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78,-181.5,-70.5,-181.5</points>
<connection>
<GID>213</GID>
<name>IN_4</name></connection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77,-184.5,-77,-182.5</points>
<intersection>-184.5 2</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77,-182.5,-70.5,-182.5</points>
<connection>
<GID>213</GID>
<name>IN_3</name></connection>
<intersection>-77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-184.5,-77,-184.5</points>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-77 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83.5,-186.5,-76,-186.5</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-76 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-76,-186.5,-76,-183.5</points>
<intersection>-186.5 1</intersection>
<intersection>-183.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-76,-183.5,-70.5,-183.5</points>
<connection>
<GID>213</GID>
<name>IN_2</name></connection>
<intersection>-76 3</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,-190.5,-74,-185.5</points>
<intersection>-190.5 2</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,-185.5,-70.5,-185.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-83.5,-190.5,-74,-190.5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>-74 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-188.5,-75,-184.5</points>
<intersection>-188.5 1</intersection>
<intersection>-184.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-83.5,-188.5,-75,-188.5</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,-184.5,-70.5,-184.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,-176.5,-67.5,-176.5</points>
<connection>
<GID>213</GID>
<name>load</name></connection>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,-214.5,-77.5,-214</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-214 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-78,-214,-77.5,-214</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71.5,-203,-71.5,-195.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>242,-259,356,-259</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>242 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>242,-262.5,242,-259</points>
<intersection>-262.5 7</intersection>
<intersection>-259 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>236.5,-262.5,242,-262.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>242 6</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-60.5,-235,-60.5,-229</points>
<intersection>-235 7</intersection>
<intersection>-229 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-62,-229,-60,-229</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>-60.5 1</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-60.5,-235,-60,-235</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>-60.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>155,-280.5,156,-280.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<connection>
<GID>262</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>158,-280.5,159,-280.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,-202,-81,-161.5</points>
<intersection>-202 10</intersection>
<intersection>-199 5</intersection>
<intersection>-195.5 13</intersection>
<intersection>-161.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-84,-161.5,-81,-161.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-81,-199,-60,-199</points>
<intersection>-81 0</intersection>
<intersection>-60 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-60,-227,-60,-199</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>-199 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-81,-202,-77.5,-202</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-83,-195.5,-81,-195.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,-196.5,-89,-196.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-286,152.5,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-286,155.5,-286</points>
<intersection>152.5 0</intersection>
<intersection>155.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152.5,-274.5,154,-274.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>152.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>155.5,-288.5,155.5,-286</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>164,-280.5,165,-280.5</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<connection>
<GID>268</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>167,-280.5,168,-280.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-286,161.5,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-286,164.5,-286</points>
<intersection>161.5 0</intersection>
<intersection>164.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161.5,-274.5,163,-274.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>161.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>164.5,-288.5,164.5,-286</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>173,-280.5,174,-280.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<connection>
<GID>272</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>176,-280.5,177,-280.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>273</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-286,170.5,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,-286,173.5,-286</points>
<intersection>170.5 0</intersection>
<intersection>173.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-274.5,172,-274.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>170.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>173.5,-288.5,173.5,-286</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>182.5,-280.5,183.5,-280.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<connection>
<GID>276</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>185.5,-280.5,186.5,-280.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>277</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-286,180,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180,-286,183,-286</points>
<intersection>180 0</intersection>
<intersection>183 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180,-274.5,181.5,-274.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>180 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>183,-288.5,183,-286</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>191.5,-280.5,192.5,-280.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<connection>
<GID>280</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>194.5,-280.5,195.5,-280.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-286,189,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-286,192,-286</points>
<intersection>189 0</intersection>
<intersection>192 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189,-274.5,190.5,-274.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>189 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>192,-288.5,192,-286</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>200.5,-280.5,201.5,-280.5</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<connection>
<GID>284</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>203.5,-280.5,204.5,-280.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<connection>
<GID>285</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-286,198,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-286,201,-286</points>
<intersection>198 0</intersection>
<intersection>201 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-274.5,199.5,-274.5</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201,-288.5,201,-286</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>209.5,-280.5,210.5,-280.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<connection>
<GID>288</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>212.5,-280.5,213.5,-280.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<connection>
<GID>289</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-286,207,-274.5</points>
<intersection>-286 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-286,210,-286</points>
<intersection>207 0</intersection>
<intersection>210 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>207,-274.5,208.5,-274.5</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>210,-288.5,210,-286</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>-286 1</intersection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-74,-226.5,-68,-226.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>-68 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-68,-230,-68,-226.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-226.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-213.5,-57,-206</points>
<intersection>-213.5 1</intersection>
<intersection>-206 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,-213.5,7,-213.5</points>
<intersection>-57 0</intersection>
<intersection>-54 3</intersection>
<intersection>-47.5 10</intersection>
<intersection>-38.5 9</intersection>
<intersection>-29 8</intersection>
<intersection>-20 7</intersection>
<intersection>-11 6</intersection>
<intersection>-2 5</intersection>
<intersection>7 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-206,-56.5,-206</points>
<connection>
<GID>179</GID>
<name>clock</name></connection>
<intersection>-57 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-54,-228,-54,-213.5</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>7,-244.5,7,-206</points>
<connection>
<GID>212</GID>
<name>clock</name></connection>
<intersection>-244.5 12</intersection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-2,-213.5,-2,-206</points>
<connection>
<GID>208</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-11,-213.5,-11,-206</points>
<connection>
<GID>204</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-20,-213.5,-20,-206</points>
<connection>
<GID>200</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-29,-213.5,-29,-206</points>
<connection>
<GID>196</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-38.5,-213.5,-38.5,-206</points>
<connection>
<GID>192</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-47.5,-213.5,-47.5,-206</points>
<connection>
<GID>187</GID>
<name>clock</name></connection>
<intersection>-213.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>7,-244.5,92.5,-244.5</points>
<intersection>7 4</intersection>
<intersection>92.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>92.5,-320,92.5,-182</points>
<intersection>-320 24</intersection>
<intersection>-311.5 31</intersection>
<intersection>-303 30</intersection>
<intersection>-295 29</intersection>
<intersection>-287.5 28</intersection>
<intersection>-280 27</intersection>
<intersection>-272.5 26</intersection>
<intersection>-265 25</intersection>
<intersection>-244.5 12</intersection>
<intersection>-237 16</intersection>
<intersection>-228.5 22</intersection>
<intersection>-220 21</intersection>
<intersection>-212 20</intersection>
<intersection>-204.5 19</intersection>
<intersection>-197 18</intersection>
<intersection>-189.5 17</intersection>
<intersection>-182 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>87.5,-182,92.5,-182</points>
<connection>
<GID>228</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>87.5,-237,112.5,-237</points>
<connection>
<GID>221</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection>
<intersection>112.5 35</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>87.5,-189.5,92.5,-189.5</points>
<connection>
<GID>227</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>87.5,-197,92.5,-197</points>
<connection>
<GID>226</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>87.5,-204.5,92.5,-204.5</points>
<connection>
<GID>225</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>87.5,-212,92.5,-212</points>
<connection>
<GID>224</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>87.5,-220,92.5,-220</points>
<connection>
<GID>223</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>87.5,-228.5,92.5,-228.5</points>
<connection>
<GID>222</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>89.5,-320,114.5,-320</points>
<connection>
<GID>231</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection>
<intersection>114.5 33</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>89.5,-265,92.5,-265</points>
<connection>
<GID>238</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>89.5,-272.5,92.5,-272.5</points>
<connection>
<GID>237</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>89.5,-280,92.5,-280</points>
<connection>
<GID>236</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>89.5,-287.5,92.5,-287.5</points>
<connection>
<GID>235</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>89.5,-295,92.5,-295</points>
<connection>
<GID>234</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>89.5,-303,92.5,-303</points>
<connection>
<GID>233</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>89.5,-311.5,92.5,-311.5</points>
<connection>
<GID>232</GID>
<name>clock</name></connection>
<intersection>92.5 13</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>114.5,-320,114.5,-300</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-320 24</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>112.5,-237,112.5,-217</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-237 16</intersection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-288.5,157,-286.5</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-288.5,158.5,-288.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-288.5,175,-286.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-288.5,177,-288.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-288.5,166,-286.5</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-288.5,167.5,-288.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-288.5,184.5,-286.5</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-288.5,186,-288.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-288.5,193.5,-286.5</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-288.5,195,-288.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202.5,-288.5,202.5,-286.5</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202.5,-288.5,204,-288.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>202.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211.5,-288.5,211.5,-286.5</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211.5,-288.5,213,-288.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-223.5,-34,-219</points>
<intersection>-223.5 16</intersection>
<intersection>-222.5 8</intersection>
<intersection>-221.5 7</intersection>
<intersection>-219 18</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-34,-221.5,-33,-221.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-34.5,-222.5,-34,-222.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-34,-223.5,-33,-223.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-34,-219,-33,-219</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-94,-216,-94,-216</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54.5,-188.5,8.5,-188.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>-46 4</intersection>
<intersection>-37 6</intersection>
<intersection>-28 7</intersection>
<intersection>-18.5 8</intersection>
<intersection>-9.5 9</intersection>
<intersection>-0.5 10</intersection>
<intersection>8.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8.5,-189,8.5,-188.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-46,-189,-46,-188.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-37,-189,-37,-188.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-28,-189,-28,-188.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-18.5,-189,-18.5,-188.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-9.5,-189,-9.5,-188.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-0.5,-189,-0.5,-188.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-188.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-44.5,-222.5,-38.5,-222.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<connection>
<GID>266</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,-189,-50,-187</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,-187,4.5,-187</points>
<intersection>-60.5 2</intersection>
<intersection>-50 0</intersection>
<intersection>-41 5</intersection>
<intersection>-32 6</intersection>
<intersection>-22.5 7</intersection>
<intersection>-13.5 8</intersection>
<intersection>-4.5 9</intersection>
<intersection>4.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-60.5,-194.5,-60.5,-187</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>4.5,-189,4.5,-187</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-41,-189,-41,-187</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-32,-189,-32,-187</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-22.5,-189,-22.5,-187</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-13.5,-189,-13.5,-187</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-4.5,-189,-4.5,-187</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-187 1</intersection></vsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-70.5,-187.5,-67.5,-187.5</points>
<connection>
<GID>292</GID>
<name>CLK</name></connection>
<connection>
<GID>213</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>153.5,-221,154.5,-221</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<connection>
<GID>295</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>156.5,-221,157.5,-221</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>236,-322,238.5,-322</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>236 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>236,-323.5,236,-322</points>
<intersection>-323.5 12</intersection>
<intersection>-322 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>230,-323.5,236,-323.5</points>
<connection>
<GID>331</GID>
<name>CLK</name></connection>
<intersection>236 11</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-318,232,-318</points>
<connection>
<GID>335</GID>
<name>OUT_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-226.5,151,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-226.5,154,-226.5</points>
<intersection>151 0</intersection>
<intersection>154 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-215,152.5,-215</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>154,-229,154,-226.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>162.5,-221,163.5,-221</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<connection>
<GID>304</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>165.5,-221,166.5,-221</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<connection>
<GID>305</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-226.5,160,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-226.5,163,-226.5</points>
<intersection>160 0</intersection>
<intersection>163 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-215,161.5,-215</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>163,-229,163,-226.5</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>171.5,-221,172.5,-221</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<connection>
<GID>308</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>174.5,-221,175.5,-221</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>309</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-226.5,169,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169,-226.5,172,-226.5</points>
<intersection>169 0</intersection>
<intersection>172 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-215,170.5,-215</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>169 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>172,-229,172,-226.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>181,-221,182,-221</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<connection>
<GID>312</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,-221,185,-221</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-226.5,178.5,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-226.5,181.5,-226.5</points>
<intersection>178.5 0</intersection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-215,180,-215</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>178.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>181.5,-229,181.5,-226.5</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>190,-221,191,-221</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<connection>
<GID>316</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>193,-221,194,-221</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<connection>
<GID>317</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-226.5,187.5,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,-226.5,190.5,-226.5</points>
<intersection>187.5 0</intersection>
<intersection>190.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-215,189,-215</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>190.5,-229,190.5,-226.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>199,-221,200,-221</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<connection>
<GID>320</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>202,-221,203,-221</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<connection>
<GID>321</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-226.5,196.5,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,-226.5,199.5,-226.5</points>
<intersection>196.5 0</intersection>
<intersection>199.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196.5,-215,198,-215</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>196.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>199.5,-229,199.5,-226.5</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>208,-221,209,-221</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<connection>
<GID>324</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>211,-221,212,-221</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>325</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205.5,-226.5,205.5,-215</points>
<intersection>-226.5 1</intersection>
<intersection>-215 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205.5,-226.5,208.5,-226.5</points>
<intersection>205.5 0</intersection>
<intersection>208.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>205.5,-215,207,-215</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>205.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>208.5,-229,208.5,-226.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238.5,-320,238.5,-319</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>-319 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>238,-319,238.5,-319</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>238.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>224.5,-320,232,-320</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>224.5 14</intersection>
<intersection>230.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>230.5,-325.5,230.5,-320</points>
<intersection>-325.5 16</intersection>
<intersection>-320 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>224.5,-320,224.5,-314.5</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>-320 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>230.5,-325.5,237,-325.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>230.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-229,155.5,-227</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-229,157,-229</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-229,173.5,-227</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,-229,175.5,-229</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-229,164.5,-227</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164.5,-229,166,-229</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-229,183,-227</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-229,184.5,-229</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-229,192,-227</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-229,193.5,-229</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-229,201,-227</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,-229,202.5,-229</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-229,210,-227</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210,-229,211.5,-229</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-325.5,248,-321</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>-325.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>241,-325.5,248,-325.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-314,247,-314</points>
<connection>
<GID>333</GID>
<name>clock</name></connection>
<intersection>247 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>247,-315,247,-314</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>-314 1</intersection></vsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,-195.5,-66.5,-188.5</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-195.5 8</intersection>
<intersection>-188.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-66.5,-188.5,-58.5,-188.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-67.5,-195.5,-66.5,-195.5</points>
<connection>
<GID>403</GID>
<name>OUT_0</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-313,235,-313</points>
<connection>
<GID>333</GID>
<name>count_enable</name></connection>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228,-318,228,-302</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>-302 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228,-302,244,-302</points>
<intersection>228 0</intersection>
<intersection>239.5 3</intersection>
<intersection>244 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>244,-312,244,-302</points>
<connection>
<GID>333</GID>
<name>clear</name></connection>
<intersection>-302 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>239.5,-302.5,239.5,-302</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>-302 1</intersection></vsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>238,-309,238,-308.5</points>
<connection>
<GID>333</GID>
<name>OUT_3</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>238,-308.5,238.5,-308.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>238 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241,-309,241,-308.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>-308.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>240.5,-308.5,241,-308.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>241 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>238,-298.5,247,-298.5</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>244.5,-322,251.5,-322</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>244.5 35</intersection>
<intersection>246 34</intersection>
<intersection>251.5 37</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>246,-322,246,-321</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-322 6</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>244.5,-322,244.5,-321</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>-322 6</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>251.5,-322,251.5,-320</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-322 6</intersection></vsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>224.5,-310.5,224.5,-310.5</points>
<connection>
<GID>303</GID>
<name>OUT_0</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-298.5,251,-294.5</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-294.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>251,-294.5,258.5,-294.5</points>
<intersection>251 0</intersection>
<intersection>258.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>258.5,-294.5,258.5,-290.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>-294.5 27</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>224.5,-306.5,224.5,-295.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>-299.5 10</intersection>
<intersection>-295.5 43</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>224.5,-299.5,228,-299.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>224.5 7</intersection>
<intersection>228 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>228,-299.5,228,-297.5</points>
<intersection>-299.5 10</intersection>
<intersection>-297.5 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>228,-297.5,232,-297.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>228 28</intersection></hsegment>
<hsegment>
<ID>43</ID>
<points>224.5,-295.5,229,-295.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>224.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232,-299.5,232,-299.5</points>
<connection>
<GID>367</GID>
<name>OUT_0</name></connection>
<connection>
<GID>390</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229,-291.5,229,-291.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>257.5,-312.5,363.5,-312.5</points>
<intersection>257.5 20</intersection>
<intersection>263 9</intersection>
<intersection>272 8</intersection>
<intersection>281 7</intersection>
<intersection>290.5 6</intersection>
<intersection>299.5 16</intersection>
<intersection>308.5 12</intersection>
<intersection>317.5 14</intersection>
<intersection>326.5 11</intersection>
<intersection>363.5 18</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>290.5,-312.5,290.5,-308.5</points>
<connection>
<GID>350</GID>
<name>clock</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>281,-312.5,281,-308.5</points>
<connection>
<GID>346</GID>
<name>clock</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>272,-312.5,272,-308.5</points>
<connection>
<GID>342</GID>
<name>clock</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>263,-312.5,263,-308.5</points>
<connection>
<GID>337</GID>
<name>clock</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>326.5,-312.5,326.5,-308.5</points>
<intersection>-312.5 2</intersection>
<intersection>-308.5 33</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>308.5,-312.5,308.5,-308.5</points>
<intersection>-312.5 2</intersection>
<intersection>-308.5 31</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>317.5,-312.5,317.5,-308.5</points>
<intersection>-312.5 2</intersection>
<intersection>-308.5 32</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>299.5,-312.5,299.5,-308.5</points>
<intersection>-312.5 2</intersection>
<intersection>-308.5 30</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>363.5,-312.5,363.5,-305.5</points>
<intersection>-312.5 2</intersection>
<intersection>-305.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>363.5,-305.5,365.5,-305.5</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>363.5 18</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>257.5,-321,257.5,-312.5</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-312.5 2</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>299,-308.5,299.5,-308.5</points>
<connection>
<GID>354</GID>
<name>clock</name></connection>
<intersection>299.5 16</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>308,-308.5,308.5,-308.5</points>
<connection>
<GID>358</GID>
<name>clock</name></connection>
<intersection>308.5 12</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>317,-308.5,317.5,-308.5</points>
<connection>
<GID>362</GID>
<name>clock</name></connection>
<intersection>317.5 14</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>326,-308.5,326.5,-308.5</points>
<connection>
<GID>366</GID>
<name>clock</name></connection>
<intersection>326.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>268.5,-297.5,269.5,-297.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<connection>
<GID>338</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>271.5,-297.5,272.5,-297.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<connection>
<GID>339</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257,-289,323.5,-289</points>
<intersection>257 27</intersection>
<intersection>269.5 42</intersection>
<intersection>278.5 34</intersection>
<intersection>287.5 37</intersection>
<intersection>296.5 38</intersection>
<intersection>305.5 39</intersection>
<intersection>314.5 40</intersection>
<intersection>323.5 36</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>257,-297.5,257,-289</points>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>278.5,-291.5,278.5,-289</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>323.5,-291.5,323.5,-289</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>287.5,-291.5,287.5,-289</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>296.5,-291.5,296.5,-289</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>305.5,-291.5,305.5,-289</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>314.5,-291.5,314.5,-289</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>269.5,-291.5,269.5,-289</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-289 1</intersection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-303,266,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-303,269,-303</points>
<intersection>266 0</intersection>
<intersection>269 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266,-291.5,267.5,-291.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>266 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>269,-305.5,269,-303</points>
<connection>
<GID>337</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>277.5,-297.5,278.5,-297.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<connection>
<GID>343</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>280.5,-297.5,281.5,-297.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>344</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-303,275,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275,-303,278,-303</points>
<intersection>275 0</intersection>
<intersection>278 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>275,-291.5,276.5,-291.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>278,-305.5,278,-303</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>286.5,-297.5,287.5,-297.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<connection>
<GID>347</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>289.5,-297.5,290.5,-297.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<connection>
<GID>348</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>284,-303,284,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284,-303,287,-303</points>
<intersection>284 0</intersection>
<intersection>287 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>284,-291.5,285.5,-291.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>284 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>287,-305.5,287,-303</points>
<connection>
<GID>346</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>295.5,-297.5,296.5,-297.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<connection>
<GID>351</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>298.5,-297.5,299.5,-297.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>352</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-303,293,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-303,296.5,-303</points>
<intersection>293 0</intersection>
<intersection>296.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>293,-291.5,294.5,-291.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>293 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>296.5,-305.5,296.5,-303</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>304.5,-297.5,305.5,-297.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<connection>
<GID>355</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>307.5,-297.5,308.5,-297.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<connection>
<GID>356</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302,-303,302,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302,-303,305,-303</points>
<intersection>302 0</intersection>
<intersection>305 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>302,-291.5,303.5,-291.5</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>302 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305,-305.5,305,-303</points>
<connection>
<GID>354</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>313.5,-297.5,314.5,-297.5</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<connection>
<GID>359</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>316.5,-297.5,317.5,-297.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<connection>
<GID>360</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-303,311,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-303,314,-303</points>
<intersection>311 0</intersection>
<intersection>314 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>311,-291.5,312.5,-291.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>311 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>314,-305.5,314,-303</points>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>322.5,-297.5,323.5,-297.5</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<connection>
<GID>363</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>325.5,-297.5,326.5,-297.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-303,320,-291.5</points>
<intersection>-303 1</intersection>
<intersection>-291.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-303,323,-303</points>
<intersection>320 0</intersection>
<intersection>323 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>320,-291.5,321.5,-291.5</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>320 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>323,-305.5,323,-303</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>-303 1</intersection></vsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-305.5,263,-288</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>-288 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>257,-288,263,-288</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<intersection>263 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-305.5,270.5,-303.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-305.5,272,-305.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288.5,-305.5,288.5,-303.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288.5,-305.5,290.5,-305.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>288.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279.5,-305.5,279.5,-303.5</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279.5,-305.5,281,-305.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>279.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297.5,-305.5,297.5,-303.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297.5,-305.5,299,-305.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>297.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>306.5,-305.5,306.5,-303.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>306.5,-305.5,308,-305.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>306.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>315.5,-305.5,315.5,-303.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>315.5,-305.5,317,-305.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>315.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>324.5,-305.5,324.5,-303.5</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>324.5,-305.5,326,-305.5</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>324.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325.5,-291.5,325.5,-281</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>-281 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-281,325.5,-281</points>
<connection>
<GID>368</GID>
<name>OUT_7</name></connection>
<intersection>325.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-291.5,316.5,-282</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>-282 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-282,316.5,-282</points>
<connection>
<GID>368</GID>
<name>OUT_6</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,-291.5,307.5,-283</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<intersection>-283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-283,307.5,-283</points>
<connection>
<GID>368</GID>
<name>OUT_5</name></connection>
<intersection>307.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>298.5,-291.5,298.5,-284</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>-284 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-284,298.5,-284</points>
<connection>
<GID>368</GID>
<name>OUT_4</name></connection>
<intersection>298.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>289.5,-291.5,289.5,-285</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-285 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-285,289.5,-285</points>
<connection>
<GID>368</GID>
<name>OUT_3</name></connection>
<intersection>289.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280.5,-291.5,280.5,-286</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-286,280.5,-286</points>
<connection>
<GID>368</GID>
<name>OUT_2</name></connection>
<intersection>280.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>252,-290,252,-290</points>
<connection>
<GID>368</GID>
<name>clock</name></connection>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-291.5,248,-288</points>
<intersection>-291.5 2</intersection>
<intersection>-288 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,-288,249,-288</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243,-291.5,248,-291.5</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-289.5,246.5,-287</points>
<intersection>-289.5 1</intersection>
<intersection>-287 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-289.5,246.5,-289.5</points>
<connection>
<GID>377</GID>
<name>OUT_0</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>246.5,-287,249,-287</points>
<connection>
<GID>368</GID>
<name>IN_1</name></connection>
<intersection>246.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-287.5,246,-286</points>
<intersection>-287.5 2</intersection>
<intersection>-286 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246,-286,249,-286</points>
<connection>
<GID>368</GID>
<name>IN_2</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243,-287.5,246,-287.5</points>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-285.5,245,-285</points>
<intersection>-285.5 1</intersection>
<intersection>-285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-285.5,245,-285.5</points>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>245,-285,249,-285</points>
<connection>
<GID>368</GID>
<name>IN_3</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-284,245,-283.5</points>
<intersection>-284 1</intersection>
<intersection>-283.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-284,249,-284</points>
<connection>
<GID>368</GID>
<name>IN_4</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243,-283.5,245,-283.5</points>
<connection>
<GID>374</GID>
<name>OUT_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,-282,247,-279.5</points>
<intersection>-282 1</intersection>
<intersection>-279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,-282,249,-282</points>
<connection>
<GID>368</GID>
<name>IN_6</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243,-279.5,247,-279.5</points>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-283,246,-281.5</points>
<intersection>-283 2</intersection>
<intersection>-281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-281.5,246,-281.5</points>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>246,-283,249,-283</points>
<connection>
<GID>368</GID>
<name>IN_5</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,-281,248,-277.5</points>
<intersection>-281 2</intersection>
<intersection>-277.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243,-277.5,248,-277.5</points>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>248,-281,249,-281</points>
<connection>
<GID>368</GID>
<name>IN_7</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>252,-279,252,-279</points>
<connection>
<GID>368</GID>
<name>load</name></connection>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-285,372,-282</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-285 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-285,372,-285</points>
<intersection>360 2</intersection>
<intersection>372 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>360,-285,360,-260</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>-285 1</intersection></vsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-276,372,-274</points>
<connection>
<GID>380</GID>
<name>OUT_0</name></connection>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-275 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372,-275,383,-275</points>
<intersection>372 0</intersection>
<intersection>383 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>383,-275,383,-254</points>
<intersection>-275 3</intersection>
<intersection>-254 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>383,-254,384,-254</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>383 4</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-268,372,-266</points>
<connection>
<GID>381</GID>
<name>OUT_0</name></connection>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-267 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372,-267,382,-267</points>
<intersection>372 0</intersection>
<intersection>382 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>382,-267,382,-253</points>
<intersection>-267 3</intersection>
<intersection>-253 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>382,-253,384,-253</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>382 4</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-260,372,-258</points>
<connection>
<GID>382</GID>
<name>OUT_0</name></connection>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>-259 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>372,-259,381,-259</points>
<intersection>372 0</intersection>
<intersection>381 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>381,-259,381,-252</points>
<intersection>-259 6</intersection>
<intersection>-252 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>381,-252,384,-252</points>
<connection>
<GID>379</GID>
<name>IN_2</name></connection>
<intersection>381 7</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-252,372,-250</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>-251 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372,-251,384,-251</points>
<connection>
<GID>379</GID>
<name>IN_3</name></connection>
<intersection>372 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-250,380,-243</points>
<intersection>-250 5</intersection>
<intersection>-243 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>380,-250,384,-250</points>
<connection>
<GID>379</GID>
<name>IN_4</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>372,-243,380,-243</points>
<intersection>372 8</intersection>
<intersection>380 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>372,-244,372,-242</points>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>-243 6</intersection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-236,372,-234</points>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-235 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372,-235,381,-235</points>
<intersection>372 0</intersection>
<intersection>381 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>381,-249,381,-235</points>
<intersection>-249 5</intersection>
<intersection>-235 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>381,-249,384,-249</points>
<connection>
<GID>379</GID>
<name>IN_5</name></connection>
<intersection>381 4</intersection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-228,372,-226</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-227 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>372,-227,382,-227</points>
<intersection>372 0</intersection>
<intersection>382 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>382,-248,382,-227</points>
<intersection>-248 5</intersection>
<intersection>-227 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>382,-248,384,-248</points>
<connection>
<GID>379</GID>
<name>IN_6</name></connection>
<intersection>382 4</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>372,-220,372,-219</points>
<connection>
<GID>387</GID>
<name>OUT_0</name></connection>
<intersection>-219 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>372,-219,383,-219</points>
<intersection>372 0</intersection>
<intersection>383 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>383,-247,383,-219</points>
<intersection>-247 3</intersection>
<intersection>-219 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>383,-247,384,-247</points>
<connection>
<GID>379</GID>
<name>IN_7</name></connection>
<intersection>383 2</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>387,-245,387,-245</points>
<connection>
<GID>379</GID>
<name>load</name></connection>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344,-305.5,344,-261</points>
<intersection>-305.5 2</intersection>
<intersection>-261 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,-261,356,-261</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>344 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>332,-305.5,344,-305.5</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<intersection>344 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-291.5,273.5,-290.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262.5,-290.5,327.5,-290.5</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>273.5 0</intersection>
<intersection>282.5 5</intersection>
<intersection>291.5 6</intersection>
<intersection>300.5 7</intersection>
<intersection>309.5 8</intersection>
<intersection>318.5 9</intersection>
<intersection>327.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>327.5,-291.5,327.5,-290.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>282.5,-291.5,282.5,-290.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>291.5,-291.5,291.5,-290.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>300.5,-291.5,300.5,-290.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>309.5,-291.5,309.5,-290.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>318.5,-291.5,318.5,-290.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-290.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229,-287.5,233,-287.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<connection>
<GID>399</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212.5,-274.5,212.5,-263.5</points>
<connection>
<GID>289</GID>
<name>IN_1</name></connection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-263.5,212.5,-263.5</points>
<intersection>130.5 2</intersection>
<intersection>212.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>130.5,-287,130.5,-263.5</points>
<intersection>-287 3</intersection>
<intersection>-263.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-287,130.5,-287</points>
<connection>
<GID>230</GID>
<name>OUT_7</name></connection>
<intersection>130.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-229,136.5,-211</points>
<intersection>-229 1</intersection>
<intersection>-211 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-229,148,-229</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117.5,-211,136.5,-211</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-215,156.5,-210</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-210,156.5,-210</points>
<connection>
<GID>220</GID>
<name>OUT_1</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>165.5,-215,165.5,-209</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>-209 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-209,165.5,-209</points>
<connection>
<GID>220</GID>
<name>OUT_2</name></connection>
<intersection>165.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-215,174.5,-208</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-208,174.5,-208</points>
<connection>
<GID>220</GID>
<name>OUT_3</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-215,184,-207</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-207,184,-207</points>
<connection>
<GID>220</GID>
<name>OUT_4</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>386</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>144.5,-273,144.5,-173</points>
<intersection>-273 59</intersection>
<intersection>-213 37</intersection>
<intersection>-173 35</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>17.5,-222.5,17.5,-173</points>
<intersection>-222.5 88</intersection>
<intersection>-173 35</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>17.5,-173,144.5,-173</points>
<intersection>17.5 22</intersection>
<intersection>144.5 2</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>144.5,-213,209,-213</points>
<intersection>144.5 2</intersection>
<intersection>154.5 80</intersection>
<intersection>163.5 52</intersection>
<intersection>172.5 53</intersection>
<intersection>182 54</intersection>
<intersection>191 55</intersection>
<intersection>200 56</intersection>
<intersection>209 51</intersection></hsegment>
<vsegment>
<ID>51</ID>
<points>209,-215,209,-213</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>163.5,-215,163.5,-213</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>172.5,-215,172.5,-213</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>182,-215,182,-213</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>191,-215,191,-213</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>200,-215,200,-213</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<hsegment>
<ID>59</ID>
<points>144.5,-273,210.5,-273</points>
<intersection>144.5 2</intersection>
<intersection>156 60</intersection>
<intersection>165 74</intersection>
<intersection>174 75</intersection>
<intersection>183.5 76</intersection>
<intersection>192.5 77</intersection>
<intersection>201.5 78</intersection>
<intersection>210.5 73</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>156,-274.5,156,-273</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>210.5,-274.5,210.5,-273</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>165,-274.5,165,-273</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>174,-274.5,174,-273</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>183.5,-274.5,183.5,-273</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>192.5,-274.5,192.5,-273</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>201.5,-274.5,201.5,-273</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-273 59</intersection></vsegment>
<vsegment>
<ID>80</ID>
<points>154.5,-215,154.5,-213</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>-213 37</intersection></vsegment>
<hsegment>
<ID>88</ID>
<points>-27,-222.5,17.5,-222.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<intersection>17.5 22</intersection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202,-215,202,-205</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>-205 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-205,202,-205</points>
<connection>
<GID>220</GID>
<name>OUT_6</name></connection>
<intersection>202 0</intersection></hsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-215,211,-204</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>-204 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-204,211,-204</points>
<connection>
<GID>220</GID>
<name>OUT_7</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-294,137.5,-288.5</points>
<intersection>-294 1</intersection>
<intersection>-288.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-294,137.5,-294</points>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-288.5,149.5,-288.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-274.5,158,-269.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>-269.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-269.5,158,-269.5</points>
<intersection>136.5 2</intersection>
<intersection>158 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>136.5,-293,136.5,-269.5</points>
<intersection>-293 5</intersection>
<intersection>-269.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>119.5,-293,136.5,-293</points>
<connection>
<GID>230</GID>
<name>OUT_1</name></connection>
<intersection>136.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-274.5,167,-268.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-268.5,167,-268.5</points>
<intersection>135.5 2</intersection>
<intersection>167 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>135.5,-292,135.5,-268.5</points>
<intersection>-292 3</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-292,135.5,-292</points>
<connection>
<GID>230</GID>
<name>OUT_2</name></connection>
<intersection>135.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-274.5,176,-267.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>-267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-267.5,176,-267.5</points>
<intersection>134.5 2</intersection>
<intersection>176 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>134.5,-291,134.5,-267.5</points>
<intersection>-291 3</intersection>
<intersection>-267.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-291,134.5,-291</points>
<connection>
<GID>230</GID>
<name>OUT_3</name></connection>
<intersection>134.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-274.5,185.5,-266.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>-266.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-266.5,185.5,-266.5</points>
<intersection>133.5 2</intersection>
<intersection>185.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>133.5,-290,133.5,-266.5</points>
<intersection>-290 3</intersection>
<intersection>-266.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-290,133.5,-290</points>
<connection>
<GID>230</GID>
<name>OUT_4</name></connection>
<intersection>133.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-274.5,194.5,-265.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>-265.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,-265.5,194.5,-265.5</points>
<intersection>132.5 2</intersection>
<intersection>194.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>132.5,-289,132.5,-265.5</points>
<intersection>-289 5</intersection>
<intersection>-265.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>119.5,-289,132.5,-289</points>
<connection>
<GID>230</GID>
<name>OUT_5</name></connection>
<intersection>132.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203.5,-274.5,203.5,-264.5</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>-264.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,-264.5,203.5,-264.5</points>
<intersection>131.5 2</intersection>
<intersection>203.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>131.5,-288,131.5,-264.5</points>
<intersection>-288 3</intersection>
<intersection>-264.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>119.5,-288,131.5,-288</points>
<connection>
<GID>230</GID>
<name>OUT_6</name></connection>
<intersection>131.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379,-304.5,379,-226</points>
<intersection>-304.5 1</intersection>
<intersection>-282 4</intersection>
<intersection>-274 3</intersection>
<intersection>-266 10</intersection>
<intersection>-258 9</intersection>
<intersection>-250 8</intersection>
<intersection>-242 11</intersection>
<intersection>-234 12</intersection>
<intersection>-226 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>371.5,-304.5,387,-304.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>379 0</intersection>
<intersection>387 14</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>375,-274,379,-274</points>
<connection>
<GID>381</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>375,-282,379,-282</points>
<connection>
<GID>380</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>375,-250,379,-250</points>
<connection>
<GID>384</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>375,-258,379,-258</points>
<connection>
<GID>383</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>375,-266,379,-266</points>
<connection>
<GID>382</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>375,-242,379,-242</points>
<connection>
<GID>385</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>375,-234,379,-234</points>
<connection>
<GID>386</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>387,-304.5,387,-260</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-304.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>375,-226,379,-226</points>
<connection>
<GID>387</GID>
<name>clock</name></connection>
<intersection>379 0</intersection></hsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-291.5,271.5,-287</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>-287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-287,271.5,-287</points>
<connection>
<GID>368</GID>
<name>OUT_1</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>387,-256,387,-256</points>
<connection>
<GID>379</GID>
<name>clock</name></connection>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>-94,-212,-94,-204.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-205 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-94,-205,-90.5,-205</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>-94 7</intersection>
<intersection>-90.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>-90.5,-205,-90.5,-203</points>
<intersection>-205 10</intersection>
<intersection>-203 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>-90.5,-203,-86.5,-203</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>-90.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-86.5,-205,-86.5,-205</points>
<connection>
<GID>401</GID>
<name>OUT_0</name></connection>
<connection>
<GID>402</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94,-200.5,-94,-200.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-213,112.5,-213</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<connection>
<GID>220</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-296,114.5,-296</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>230</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-215,193,-206</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-206,193,-206</points>
<connection>
<GID>220</GID>
<name>OUT_5</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-288.5,225.5,-265</points>
<intersection>-288.5 1</intersection>
<intersection>-265 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-288.5,225.5,-288.5</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-265,230.5,-265</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>406</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-266,224,-229</points>
<intersection>-266 2</intersection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>217.5,-229,224,-229</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>224,-266,230.5,-266</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-84,-158.5,358,-158.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<intersection>-80 13</intersection>
<intersection>358 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>358,-257.5,358,-158.5</points>
<connection>
<GID>257</GID>
<name>SEL_0</name></connection>
<intersection>-242.5 23</intersection>
<intersection>-158.5 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-80,-197.5,-80,-158.5</points>
<intersection>-197.5 14</intersection>
<intersection>-158.5 7</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-83,-197.5,-61.5,-197.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>-80 13</intersection>
<intersection>-61.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-61.5,-237,-61.5,-197.5</points>
<intersection>-237 19</intersection>
<intersection>-221.5 22</intersection>
<intersection>-197.5 14</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-61.5,-237,-60,-237</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>-61.5 18</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-61.5,-221.5,-50.5,-221.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>-61.5 18</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>238.5,-242.5,358,-242.5</points>
<intersection>238.5 24</intersection>
<intersection>358 10</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>238.5,-287.5,238.5,-242.5</points>
<intersection>-287.5 31</intersection>
<intersection>-242.5 23</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>237,-287.5,238.5,-287.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>238.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,79.5,-70,80.5</points>
<intersection>79.5 1</intersection>
<intersection>80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70,79.5,-69,79.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>-70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,80.5,-70,80.5</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<intersection>-70 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,76.5,-69,76.5</points>
<connection>
<GID>406</GID>
<name>OUT_0</name></connection>
<intersection>-69 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-69,76.5,-69,77.5</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-63,78.5,-61,78.5</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,77.5,-54,82.5</points>
<intersection>77.5 2</intersection>
<intersection>82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,82.5,-53,82.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,77.5,-54,77.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-71,70.5,-69,70.5</points>
<connection>
<GID>409</GID>
<name>OUT_0</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,70.5,-62,76.5</points>
<intersection>70.5 2</intersection>
<intersection>76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,76.5,-61,76.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,70.5,-62,70.5</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,79.5,-39,82.5</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,79.5,-39,79.5</points>
<intersection>-45 3</intersection>
<intersection>-39 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-45,76.5,-45,79.5</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-47,83.5,-45,83.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-47,63.5,-45,63.5</points>
<connection>
<GID>425</GID>
<name>OUT_0</name></connection>
<connection>
<GID>426</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,61.5,-45,61.5</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<intersection>-58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-58,61.5,-58,74.5</points>
<intersection>61.5 1</intersection>
<intersection>74.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-58,74.5,-45,74.5</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<intersection>-58 3</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,78.5,-46,81.5</points>
<intersection>78.5 2</intersection>
<intersection>81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,81.5,-45,81.5</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>-46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46,78.5,-38,78.5</points>
<intersection>-46 0</intersection>
<intersection>-38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-38,75.5,-38,78.5</points>
<intersection>75.5 4</intersection>
<intersection>78.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-39,75.5,-34,75.5</points>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<intersection>-38 3</intersection>
<intersection>-37 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-37,69.5,-37,75.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>75.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,67.5,-37,67.5</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>429</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,68.5,-29,68.5</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,59.5,-34,62.5</points>
<intersection>59.5 1</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,59.5,-29,59.5</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-39,62.5,-34,62.5</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,60.5,-22,63.5</points>
<intersection>60.5 2</intersection>
<intersection>63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,63.5,-22,63.5</points>
<intersection>-30 3</intersection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23,60.5,-20,60.5</points>
<connection>
<GID>422</GID>
<name>N_in0</name></connection>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<intersection>-22 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30,63.5,-30,66.5</points>
<intersection>63.5 1</intersection>
<intersection>66.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-30,66.5,-29,66.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>-30 3</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,84.5,-53,84.5</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,64.5,-23,67.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,64.5,-23,64.5</points>
<intersection>-29 3</intersection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-29,61.5,-29,64.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-391,-58,-387</points>
<intersection>-391 29</intersection>
<intersection>-387 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,-387,-56,-387</points>
<connection>
<GID>608</GID>
<name>J</name></connection>
<connection>
<GID>610</GID>
<name>OUT_0</name></connection>
<intersection>-58 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>-58,-391,-56,-391</points>
<connection>
<GID>608</GID>
<name>K</name></connection>
<intersection>-58 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-57,-395,-15,-395</points>
<intersection>-57 23</intersection>
<intersection>-26 24</intersection>
<intersection>-15 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-15,-407,-15,-395</points>
<connection>
<GID>626</GID>
<name>carry_out</name></connection>
<intersection>-395 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-57,-395,-57,-389</points>
<intersection>-395 1</intersection>
<intersection>-389 25</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>-26,-395,-26,-389</points>
<intersection>-395 1</intersection>
<intersection>-389 26</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>-57,-389,-56,-389</points>
<connection>
<GID>608</GID>
<name>clock</name></connection>
<intersection>-57 23</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-26,-389,-25,-389</points>
<connection>
<GID>609</GID>
<name>clock</name></connection>
<intersection>-26 24</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>-44,-392,-41,-392</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<connection>
<GID>614</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-49,-390,-41,-390</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>-49 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-49,-391,-49,-390</points>
<intersection>-391 8</intersection>
<intersection>-390 5</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-50,-391,-49,-391</points>
<connection>
<GID>608</GID>
<name>nQ</name></connection>
<intersection>-49 7</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-34,-388,-33,-388</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>-34 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-34,-388,-34,-387</points>
<intersection>-388 5</intersection>
<intersection>-387 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-35,-387,-34,-387</points>
<connection>
<GID>612</GID>
<name>OUT</name></connection>
<intersection>-34 6</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-34,-390,-33,-390</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<intersection>-34 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-34,-391,-34,-390</points>
<intersection>-391 7</intersection>
<intersection>-390 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-35,-391,-34,-391</points>
<connection>
<GID>613</GID>
<name>OUT</name></connection>
<intersection>-34 6</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-391,-27,-387</points>
<connection>
<GID>615</GID>
<name>OUT</name></connection>
<intersection>-391 3</intersection>
<intersection>-387 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,-387,-25,-387</points>
<connection>
<GID>609</GID>
<name>J</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27,-391,-25,-391</points>
<connection>
<GID>609</GID>
<name>K</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-419,-18,-418</points>
<connection>
<GID>626</GID>
<name>clock</name></connection>
<intersection>-419 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-48,-419,-18,-419</points>
<intersection>-48 6</intersection>
<intersection>-18 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-48,-419,-48,-403</points>
<intersection>-419 5</intersection>
<intersection>-403 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-50,-403,-48,-403</points>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection>
<intersection>-48 6</intersection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>-18.5,-405.5,-18.5,-403</points>
<intersection>-405.5 34</intersection>
<intersection>-403 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-20,-403,-17,-403</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<intersection>-18.5 5</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>-18.5,-405.5,-18,-405.5</points>
<intersection>-18.5 5</intersection>
<intersection>-18 41</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>-18,-407,-18,-405.5</points>
<connection>
<GID>626</GID>
<name>load</name></connection>
<intersection>-405.5 34</intersection></vsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-17,-407,-17,-407</points>
<connection>
<GID>623</GID>
<name>OUT_0</name></connection>
<connection>
<GID>626</GID>
<name>count_enable</name></connection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-407,-16,-401</points>
<connection>
<GID>626</GID>
<name>count_up</name></connection>
<intersection>-401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,-401,-16,-401</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<intersection>-48 2</intersection>
<intersection>-16 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-48,-401,-48,-386</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>-401 1</intersection>
<intersection>-386 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-48,-386,-41,-386</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>-48 2</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-462.5,-4,-394.5</points>
<intersection>-462.5 3</intersection>
<intersection>-409 2</intersection>
<intersection>-394.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-394.5,-3,-394.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13,-409,-4,-409</points>
<connection>
<GID>626</GID>
<name>OUT_7</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4,-462.5,1,-462.5</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-458.5,-5,-390.5</points>
<intersection>-458.5 3</intersection>
<intersection>-410 2</intersection>
<intersection>-390.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-390.5,-3,-390.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13,-410,-5,-410</points>
<connection>
<GID>626</GID>
<name>OUT_6</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5,-458.5,1,-458.5</points>
<connection>
<GID>769</GID>
<name>IN_1</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-454.5,-6,-386.5</points>
<intersection>-454.5 4</intersection>
<intersection>-411 5</intersection>
<intersection>-386.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-386.5,-3,-386.5</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-6,-454.5,1,-454.5</points>
<connection>
<GID>768</GID>
<name>IN_1</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-13,-411,-6,-411</points>
<connection>
<GID>626</GID>
<name>OUT_5</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-450.5,-7,-382.5</points>
<intersection>-450.5 4</intersection>
<intersection>-412 2</intersection>
<intersection>-382.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-382.5,-3,-382.5</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13,-412,-7,-412</points>
<connection>
<GID>626</GID>
<name>OUT_4</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-7,-450.5,1,-450.5</points>
<connection>
<GID>767</GID>
<name>IN_1</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-446.5,-8,-378.5</points>
<intersection>-446.5 4</intersection>
<intersection>-413 1</intersection>
<intersection>-378.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-413,-8,-413</points>
<connection>
<GID>626</GID>
<name>OUT_3</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-378.5,-3,-378.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-8,-446.5,1,-446.5</points>
<connection>
<GID>766</GID>
<name>IN_1</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-442.5,-9,-374.5</points>
<intersection>-442.5 3</intersection>
<intersection>-414 1</intersection>
<intersection>-374.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-414,-9,-414</points>
<connection>
<GID>626</GID>
<name>OUT_2</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-9,-374.5,-3,-374.5</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-9,-442.5,1,-442.5</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-438.5,-10,-370.5</points>
<intersection>-438.5 3</intersection>
<intersection>-415 1</intersection>
<intersection>-370.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-415,-10,-415</points>
<connection>
<GID>626</GID>
<name>OUT_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-370.5,-3,-370.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10,-438.5,1,-438.5</points>
<connection>
<GID>764</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-434.5,-11,-366.5</points>
<intersection>-434.5 3</intersection>
<intersection>-416 1</intersection>
<intersection>-366.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-416,-11,-416</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,-366.5,-3,-366.5</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-11,-434.5,1,-434.5</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-363.5,21,-363.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>16,-399.5,16,-365.5</points>
<intersection>-399.5 19</intersection>
<intersection>-365.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-365.5,21,-365.5</points>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<connection>
<GID>753</GID>
<name>OUT</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>16,-399.5,21,-399.5</points>
<connection>
<GID>666</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-403.5,15,-369.5</points>
<intersection>-403.5 3</intersection>
<intersection>-369.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-369.5,21,-369.5</points>
<connection>
<GID>651</GID>
<name>IN_1</name></connection>
<connection>
<GID>754</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>15,-403.5,21,-403.5</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-407.5,14,-373.5</points>
<intersection>-407.5 3</intersection>
<intersection>-373.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-373.5,21,-373.5</points>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14,-407.5,21,-407.5</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>13,-411.5,13,-377.5</points>
<intersection>-411.5 5</intersection>
<intersection>-377.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>13,-411.5,21,-411.5</points>
<connection>
<GID>669</GID>
<name>IN_1</name></connection>
<intersection>13 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-377.5,21,-377.5</points>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<connection>
<GID>756</GID>
<name>OUT</name></connection>
<intersection>13 4</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>12,-415.5,12,-381.5</points>
<intersection>-415.5 4</intersection>
<intersection>-381.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12,-415.5,21,-415.5</points>
<connection>
<GID>670</GID>
<name>IN_1</name></connection>
<intersection>12 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-381.5,21,-381.5</points>
<connection>
<GID>654</GID>
<name>IN_1</name></connection>
<connection>
<GID>757</GID>
<name>OUT</name></connection>
<intersection>12 3</intersection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-385.5,21,-385.5</points>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<connection>
<GID>758</GID>
<name>OUT</name></connection>
<intersection>11 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>11,-419.5,11,-385.5</points>
<intersection>-419.5 4</intersection>
<intersection>-385.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>11,-419.5,21,-419.5</points>
<connection>
<GID>671</GID>
<name>IN_1</name></connection>
<intersection>11 3</intersection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-389.5,21,-389.5</points>
<connection>
<GID>656</GID>
<name>IN_1</name></connection>
<connection>
<GID>759</GID>
<name>OUT</name></connection>
<intersection>10 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10,-423.5,10,-389.5</points>
<intersection>-423.5 4</intersection>
<intersection>-389.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>10,-423.5,21,-423.5</points>
<connection>
<GID>672</GID>
<name>IN_1</name></connection>
<intersection>10 3</intersection></hsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>9,-427.5,9,-393.5</points>
<intersection>-427.5 4</intersection>
<intersection>-393.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,-427.5,21,-427.5</points>
<connection>
<GID>673</GID>
<name>IN_1</name></connection>
<intersection>9 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>7,-393.5,21,-393.5</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<intersection>9 3</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-391.5,21,-391.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-387.5,21,-387.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<connection>
<GID>686</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-383.5,21,-383.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<connection>
<GID>685</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-379.5,21,-379.5</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<connection>
<GID>684</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-375.5,21,-375.5</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-371.5,21,-371.5</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<connection>
<GID>682</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-367.5,21,-367.5</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<connection>
<GID>681</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-431.5,21,-431.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>9,-467.5,9,-433.5</points>
<intersection>-467.5 19</intersection>
<intersection>-433.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-433.5,21,-433.5</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<connection>
<GID>763</GID>
<name>OUT</name></connection>
<intersection>9 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>9,-467.5,21,-467.5</points>
<connection>
<GID>706</GID>
<name>IN_1</name></connection>
<intersection>9 3</intersection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-471.5,10,-437.5</points>
<intersection>-471.5 3</intersection>
<intersection>-437.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-437.5,21,-437.5</points>
<connection>
<GID>691</GID>
<name>IN_1</name></connection>
<connection>
<GID>764</GID>
<name>OUT</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10,-471.5,21,-471.5</points>
<connection>
<GID>707</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-475.5,11,-441.5</points>
<intersection>-475.5 3</intersection>
<intersection>-441.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-441.5,21,-441.5</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<connection>
<GID>765</GID>
<name>OUT</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11,-475.5,21,-475.5</points>
<connection>
<GID>708</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>12,-479.5,12,-445.5</points>
<intersection>-479.5 5</intersection>
<intersection>-445.5 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>12,-479.5,21,-479.5</points>
<connection>
<GID>709</GID>
<name>IN_1</name></connection>
<intersection>12 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-445.5,21,-445.5</points>
<connection>
<GID>693</GID>
<name>IN_1</name></connection>
<connection>
<GID>766</GID>
<name>OUT</name></connection>
<intersection>12 4</intersection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>13,-483.5,13,-449.5</points>
<intersection>-483.5 4</intersection>
<intersection>-449.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13,-483.5,21,-483.5</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<intersection>13 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-449.5,21,-449.5</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<connection>
<GID>767</GID>
<name>OUT</name></connection>
<intersection>13 3</intersection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>14,-487.5,14,-453.5</points>
<intersection>-487.5 4</intersection>
<intersection>-453.5 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14,-487.5,21,-487.5</points>
<connection>
<GID>711</GID>
<name>IN_1</name></connection>
<intersection>14 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-453.5,21,-453.5</points>
<connection>
<GID>695</GID>
<name>IN_1</name></connection>
<connection>
<GID>768</GID>
<name>OUT</name></connection>
<intersection>14 3</intersection></hsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-457.5,21,-457.5</points>
<connection>
<GID>696</GID>
<name>IN_1</name></connection>
<connection>
<GID>769</GID>
<name>OUT</name></connection>
<intersection>15 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-491.5,15,-457.5</points>
<intersection>-491.5 4</intersection>
<intersection>-457.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,-491.5,21,-491.5</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>15 3</intersection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>16,-495.5,16,-461.5</points>
<intersection>-495.5 4</intersection>
<intersection>-461.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-495.5,21,-495.5</points>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>7,-461.5,21,-461.5</points>
<connection>
<GID>697</GID>
<name>IN_1</name></connection>
<connection>
<GID>770</GID>
<name>OUT</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-459.5,21,-459.5</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-493.5,8,-360</points>
<intersection>-493.5 18</intersection>
<intersection>-489.5 17</intersection>
<intersection>-485.5 16</intersection>
<intersection>-481.5 15</intersection>
<intersection>-477.5 14</intersection>
<intersection>-473.5 13</intersection>
<intersection>-469.5 12</intersection>
<intersection>-465.5 11</intersection>
<intersection>-459.5 2</intersection>
<intersection>-455.5 9</intersection>
<intersection>-451.5 8</intersection>
<intersection>-447.5 7</intersection>
<intersection>-443.5 6</intersection>
<intersection>-439.5 5</intersection>
<intersection>-435.5 4</intersection>
<intersection>-431.5 3</intersection>
<intersection>-425.5 38</intersection>
<intersection>-421.5 37</intersection>
<intersection>-417.5 36</intersection>
<intersection>-413.5 35</intersection>
<intersection>-409.5 34</intersection>
<intersection>-405.5 33</intersection>
<intersection>-401.5 32</intersection>
<intersection>-397.5 31</intersection>
<intersection>-391.5 22</intersection>
<intersection>-387.5 29</intersection>
<intersection>-383.5 28</intersection>
<intersection>-379.5 27</intersection>
<intersection>-375.5 26</intersection>
<intersection>-371.5 25</intersection>
<intersection>-367.5 24</intersection>
<intersection>-363.5 23</intersection>
<intersection>-360 21</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-459.5,17,-459.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-431.5,17,-431.5</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8,-435.5,17,-435.5</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>8,-439.5,17,-439.5</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>8,-443.5,17,-443.5</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>8,-447.5,17,-447.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8,-451.5,17,-451.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>8,-455.5,17,-455.5</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>8,-465.5,21,-465.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>8,-469.5,21,-469.5</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>8,-473.5,21,-473.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>8,-477.5,21,-477.5</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>8,-481.5,21,-481.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>8,-485.5,21,-485.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>8,-489.5,21,-489.5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>8,-493.5,21,-493.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-18,-360,8,-360</points>
<intersection>-18 40</intersection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>8,-391.5,17,-391.5</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>8,-363.5,17,-363.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>8,-367.5,17,-367.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>8,-371.5,17,-371.5</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>8,-375.5,17,-375.5</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>8,-379.5,17,-379.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>8,-383.5,17,-383.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>8,-387.5,17,-387.5</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>8,-397.5,21,-397.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>8,-401.5,21,-401.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>8,-405.5,21,-405.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>8,-409.5,21,-409.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>8,-413.5,21,-413.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>8,-417.5,21,-417.5</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>8,-421.5,21,-421.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>8,-425.5,21,-425.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>40</ID>
<points>-18,-387,-18,-360</points>
<intersection>-387 42</intersection>
<intersection>-360 21</intersection></vsegment>
<hsegment>
<ID>42</ID>
<points>-19,-387,-18,-387</points>
<connection>
<GID>609</GID>
<name>Q</name></connection>
<intersection>-18 40</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-455.5,21,-455.5</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<connection>
<GID>726</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-451.5,21,-451.5</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<connection>
<GID>725</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-447.5,21,-447.5</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<connection>
<GID>724</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-443.5,21,-443.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-439.5,21,-439.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>722</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>21,-435.5,21,-435.5</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<connection>
<GID>721</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-366.5,1,-366.5</points>
<connection>
<GID>745</GID>
<name>OUT_0</name></connection>
<connection>
<GID>753</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-370.5,1,-370.5</points>
<connection>
<GID>746</GID>
<name>OUT_0</name></connection>
<connection>
<GID>754</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-374.5,1,-374.5</points>
<connection>
<GID>747</GID>
<name>OUT_0</name></connection>
<connection>
<GID>755</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-378.5,1,-378.5</points>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection>
<connection>
<GID>756</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-382.5,1,-382.5</points>
<connection>
<GID>749</GID>
<name>OUT_0</name></connection>
<connection>
<GID>757</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-386.5,1,-386.5</points>
<connection>
<GID>750</GID>
<name>OUT_0</name></connection>
<connection>
<GID>758</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-390.5,1,-390.5</points>
<connection>
<GID>751</GID>
<name>OUT_0</name></connection>
<connection>
<GID>759</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-394.5,1,-394.5</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<connection>
<GID>760</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,-364.5,1,-364.5</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-12,-392.5,-12,-364.5</points>
<intersection>-392.5 4</intersection>
<intersection>-388.5 10</intersection>
<intersection>-384.5 9</intersection>
<intersection>-380.5 8</intersection>
<intersection>-376.5 7</intersection>
<intersection>-372.5 6</intersection>
<intersection>-368.5 5</intersection>
<intersection>-364.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12,-392.5,1,-392.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12,-368.5,1,-368.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-12,-372.5,1,-372.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-12,-376.5,1,-376.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-12,-380.5,1,-380.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-12,-384.5,1,-384.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-12,-388.5,1,-388.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-394,-12,-394</points>
<intersection>-43 12</intersection>
<intersection>-12 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-12,-460.5,-12,-394</points>
<intersection>-460.5 4</intersection>
<intersection>-456.5 10</intersection>
<intersection>-452.5 9</intersection>
<intersection>-448.5 8</intersection>
<intersection>-444.5 7</intersection>
<intersection>-440.5 6</intersection>
<intersection>-436.5 5</intersection>
<intersection>-432.5 28</intersection>
<intersection>-394 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12,-460.5,1,-460.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12,-436.5,1,-436.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-12,-440.5,1,-440.5</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-12,-444.5,1,-444.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-12,-448.5,1,-448.5</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-12,-452.5,1,-452.5</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-12,-456.5,1,-456.5</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-43,-394,-43,-364.5</points>
<intersection>-394 1</intersection>
<intersection>-388 30</intersection>
<intersection>-387 32</intersection>
<intersection>-364.5 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-43,-364.5,-17,-364.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-43 12</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-12,-432.5,1,-432.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>-43,-388,-41,-388</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<intersection>-43 12</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-50,-387,-43,-387</points>
<connection>
<GID>608</GID>
<name>Q</name></connection>
<intersection>-43 12</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39,-486,39,-486</points>
<connection>
<GID>772</GID>
<name>clock</name></connection>
<connection>
<GID>773</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>39,-475,39,-475</points>
<connection>
<GID>772</GID>
<name>load</name></connection>
<connection>
<GID>779</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-494.5,35,-477</points>
<intersection>-494.5 2</intersection>
<intersection>-477 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-477,36,-477</points>
<connection>
<GID>772</GID>
<name>IN_7</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-494.5,35,-494.5</points>
<connection>
<GID>713</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-490.5,34,-478</points>
<intersection>-490.5 2</intersection>
<intersection>-478 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-478,36,-478</points>
<connection>
<GID>772</GID>
<name>IN_6</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-490.5,34,-490.5</points>
<connection>
<GID>712</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-486.5,33,-479</points>
<intersection>-486.5 2</intersection>
<intersection>-479 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-479,36,-479</points>
<connection>
<GID>772</GID>
<name>IN_5</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-486.5,33,-486.5</points>
<connection>
<GID>711</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-482.5,32,-480</points>
<intersection>-482.5 2</intersection>
<intersection>-480 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-480,36,-480</points>
<connection>
<GID>772</GID>
<name>IN_4</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-482.5,32,-482.5</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-481,31,-478.5</points>
<intersection>-481 1</intersection>
<intersection>-478.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-481,36,-481</points>
<connection>
<GID>772</GID>
<name>IN_3</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-478.5,31,-478.5</points>
<connection>
<GID>709</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-482,30,-474.5</points>
<intersection>-482 1</intersection>
<intersection>-474.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-482,36,-482</points>
<connection>
<GID>772</GID>
<name>IN_2</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-474.5,30,-474.5</points>
<connection>
<GID>708</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-483,29,-470.5</points>
<intersection>-483 1</intersection>
<intersection>-470.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-483,36,-483</points>
<connection>
<GID>772</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-470.5,29,-470.5</points>
<connection>
<GID>707</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-484,28,-466.5</points>
<intersection>-484 1</intersection>
<intersection>-466.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-484,36,-484</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-466.5,28,-466.5</points>
<connection>
<GID>706</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>62,-435,62,-435</points>
<connection>
<GID>780</GID>
<name>clock</name></connection>
<connection>
<GID>781</GID>
<name>CLK</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 1>
<page 2>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 2>
<page 3>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 3>
<page 4>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 4>
<page 5>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 5>
<page 6>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 6>
<page 7>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 7>
<page 8>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 8>
<page 9>
<PageViewport>0,53.073,387.412,-146.734</PageViewport></page 9></circuit>