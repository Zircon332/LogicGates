<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>2.31214,-4.36478,61.1215,-65.8352</PageViewport>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>12.5,-12.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>12.5,-17.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>12.5,-22.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>17.5,-12.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>20.5,-20</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR2</type>
<position>32,-15.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>36,-15.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>12,-29</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>19,-30.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>25,-30.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-12.5,15.5,-12.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-19,16.5,-17.5</points>
<intersection>-19 3</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-17.5,16.5,-17.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16.5,-19,17.5,-19</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-22.5,16.5,-21</points>
<intersection>-22.5 2</intersection>
<intersection>-21 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-22.5,16.5,-22.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16.5,-21,17.5,-21</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-14.5,24,-12.5</points>
<intersection>-14.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-14.5,29,-14.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-12.5,24,-12.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-20,26,-16.5</points>
<intersection>-20 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-20,26,-20</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-16.5,29,-16.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-15.5,35,-15.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-29.5,15,-29</points>
<intersection>-29.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-29,15,-29</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-29.5,16,-29.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-30.5,24,-30.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 1>
<page 2>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 2>
<page 3>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 3>
<page 4>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 4>
<page 5>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 5>
<page 6>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 6>
<page 7>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 7>
<page 8>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 8>
<page 9>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 9></circuit>