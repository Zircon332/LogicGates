<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-145.91,218.771,604.184,-168.089</PageViewport>
<gate>
<ID>769</ID>
<type>AA_AND2</type>
<position>548.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>738 </input>
<output>
<ID>OUT</ID>736 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>770</ID>
<type>AA_AND2</type>
<position>552.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>748 </input>
<output>
<ID>OUT</ID>737 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1</ID>
<type>AE_FULLADDER_4BIT</type>
<position>33.5,-3</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<input>
<ID>IN_B_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<output>
<ID>OUT_1</ID>95 </output>
<output>
<ID>OUT_2</ID>96 </output>
<output>
<ID>OUT_3</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>771</ID>
<type>AE_OR2</type>
<position>550.5,-95.5</position>
<input>
<ID>IN_0</ID>737 </input>
<input>
<ID>IN_1</ID>736 </input>
<output>
<ID>OUT</ID>747 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_SMALL_INVERTER</type>
<position>7.5,7</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>772</ID>
<type>AE_DFF_LOW</type>
<position>555.5,-102.5</position>
<input>
<ID>IN_0</ID>747 </input>
<output>
<ID>OUT_0</ID>774 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>15.5,7</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>773</ID>
<type>AE_SMALL_INVERTER</type>
<position>450,-94.5</position>
<input>
<ID>IN_0</ID>712 </input>
<output>
<ID>OUT_0</ID>713 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_SMALL_INVERTER</type>
<position>23.5,7</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>774</ID>
<type>AE_REGISTER8</type>
<position>473,-80</position>
<input>
<ID>IN_0</ID>755 </input>
<input>
<ID>IN_1</ID>756 </input>
<input>
<ID>IN_2</ID>757 </input>
<input>
<ID>IN_3</ID>758 </input>
<input>
<ID>IN_4</ID>759 </input>
<input>
<ID>IN_5</ID>761 </input>
<input>
<ID>IN_6</ID>760 </input>
<input>
<ID>IN_7</ID>762 </input>
<output>
<ID>OUT_0</ID>739 </output>
<output>
<ID>OUT_1</ID>793 </output>
<output>
<ID>OUT_2</ID>753 </output>
<output>
<ID>OUT_3</ID>752 </output>
<output>
<ID>OUT_4</ID>751 </output>
<output>
<ID>OUT_5</ID>750 </output>
<output>
<ID>OUT_6</ID>749 </output>
<output>
<ID>OUT_7</ID>748 </output>
<input>
<ID>clock</ID>754 </input>
<input>
<ID>load</ID>763 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 135</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>31.5,7</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>775</ID>
<type>AA_TOGGLE</type>
<position>472,-87</position>
<output>
<ID>OUT_0</ID>754 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>38.5,3</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>776</ID>
<type>AA_TOGGLE</type>
<position>472,-72</position>
<output>
<ID>OUT_0</ID>763 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_TOGGLE</type>
<position>462,-72.5</position>
<output>
<ID>OUT_0</ID>762 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>778</ID>
<type>AA_TOGGLE</type>
<position>462,-74.5</position>
<output>
<ID>OUT_0</ID>760 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>779</ID>
<type>AA_TOGGLE</type>
<position>462,-76.5</position>
<output>
<ID>OUT_0</ID>761 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>780</ID>
<type>AA_TOGGLE</type>
<position>462,-78.5</position>
<output>
<ID>OUT_0</ID>759 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>781</ID>
<type>AA_TOGGLE</type>
<position>462,-80.5</position>
<output>
<ID>OUT_0</ID>758 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>61,40.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>782</ID>
<type>AA_TOGGLE</type>
<position>462,-82.5</position>
<output>
<ID>OUT_0</ID>757 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>783</ID>
<type>AA_TOGGLE</type>
<position>462,-84.5</position>
<output>
<ID>OUT_0</ID>756 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>784</ID>
<type>AA_TOGGLE</type>
<position>462,-86.5</position>
<output>
<ID>OUT_0</ID>755 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>785</ID>
<type>AE_REGISTER8</type>
<position>587.5,-38.5</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>766 </input>
<input>
<ID>IN_2</ID>767 </input>
<input>
<ID>IN_3</ID>768 </input>
<input>
<ID>IN_4</ID>769 </input>
<input>
<ID>IN_5</ID>770 </input>
<input>
<ID>IN_6</ID>771 </input>
<input>
<ID>IN_7</ID>772 </input>
<input>
<ID>clock</ID>794 </input>
<input>
<ID>load</ID>773 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 135</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>786</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-66.5</position>
<input>
<ID>IN_0</ID>764 </input>
<output>
<ID>OUT_0</ID>765 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>787</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-58.5</position>
<input>
<ID>IN_0</ID>765 </input>
<output>
<ID>OUT_0</ID>766 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>788</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-50.5</position>
<input>
<ID>IN_0</ID>766 </input>
<output>
<ID>OUT_0</ID>767 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>789</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-42.5</position>
<input>
<ID>IN_0</ID>767 </input>
<output>
<ID>OUT_0</ID>768 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>790</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-34.5</position>
<input>
<ID>IN_0</ID>768 </input>
<output>
<ID>OUT_0</ID>769 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>791</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-26.5</position>
<input>
<ID>IN_0</ID>769 </input>
<output>
<ID>OUT_0</ID>770 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>792</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-18.5</position>
<input>
<ID>IN_0</ID>770 </input>
<output>
<ID>OUT_0</ID>771 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>-96,52</position>
<output>
<ID>OUT_0</ID>835 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>793</ID>
<type>AE_DFF_LOW</type>
<position>573.5,-10.5</position>
<input>
<ID>IN_0</ID>771 </input>
<output>
<ID>OUT_0</ID>772 </output>
<input>
<ID>clock</ID>792 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>61,38.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>794</ID>
<type>AA_TOGGLE</type>
<position>586.5,-30.5</position>
<output>
<ID>OUT_0</ID>773 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-96,50</position>
<output>
<ID>OUT_0</ID>836 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>795</ID>
<type>AE_SMALL_INVERTER</type>
<position>586.5,-45.5</position>
<input>
<ID>IN_0</ID>792 </input>
<output>
<ID>OUT_0</ID>794 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>61,36.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>796</ID>
<type>AA_AND2</type>
<position>455,-93.5</position>
<input>
<ID>IN_0</ID>712 </input>
<input>
<ID>IN_1</ID>713 </input>
<output>
<ID>OUT</ID>706 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>-96,48</position>
<output>
<ID>OUT_0</ID>842 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>797</ID>
<type>AE_SMALL_INVERTER</type>
<position>468,-92.5</position>
<input>
<ID>IN_0</ID>706 </input>
<output>
<ID>OUT_0</ID>711 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>61,34.5</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-96,46</position>
<output>
<ID>OUT_0</ID>841 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>799</ID>
<type>AE_SMALL_INVERTER</type>
<position>480.5,-85.5</position>
<input>
<ID>IN_0</ID>711 </input>
<output>
<ID>OUT_0</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>61,22.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_AND4</type>
<position>281.5,-98.5</position>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-96,42</position>
<output>
<ID>OUT_0</ID>840 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>801</ID>
<type>AA_TOGGLE</type>
<position>123,33.5</position>
<output>
<ID>OUT_0</ID>854 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>61,20.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-96,40</position>
<output>
<ID>OUT_0</ID>839 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>803</ID>
<type>AA_TOGGLE</type>
<position>141.5,38</position>
<output>
<ID>OUT_0</ID>798 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>61,18.5</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>804</ID>
<type>AA_TOGGLE</type>
<position>141.5,40</position>
<output>
<ID>OUT_0</ID>797 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-96,38</position>
<output>
<ID>OUT_0</ID>838 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>805</ID>
<type>AA_TOGGLE</type>
<position>141.5,42</position>
<output>
<ID>OUT_0</ID>796 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>61,16.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>806</ID>
<type>AA_AND4</type>
<position>281.5,-106.5</position>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>-96,36</position>
<output>
<ID>OUT_0</ID>837 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>807</ID>
<type>AA_LABEL</type>
<position>119,33.5</position>
<gparam>LABEL_TEXT Notif</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>69,16</position>
<output>
<ID>A_greater_B</ID>26 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>103 </input>
<input>
<ID>IN_B_1</ID>104 </input>
<input>
<ID>IN_B_2</ID>105 </input>
<input>
<ID>IN_B_3</ID>106 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>808</ID>
<type>AA_LABEL</type>
<position>135,40</position>
<gparam>LABEL_TEXT Notif Index</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>809</ID>
<type>AE_SMALL_INVERTER</type>
<position>455,-82.5</position>
<input>
<ID>IN_0</ID>810 </input>
<output>
<ID>OUT_0</ID>712 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>61,4.5</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>810</ID>
<type>AE_OR2</type>
<position>567.5,-108</position>
<input>
<ID>IN_0</ID>715 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>792 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>811</ID>
<type>AE_DFF_LOW_NT</type>
<position>150.5,31.5</position>
<input>
<ID>IN_0</ID>801 </input>
<output>
<ID>OUT_0</ID>810 </output>
<input>
<ID>clock</ID>802 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>61,2.5</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>812</ID>
<type>BB_CLOCK</type>
<position>145.5,19</position>
<output>
<ID>CLK</ID>802 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>813</ID>
<type>AE_DFF_LOW_NT</type>
<position>150.5,23</position>
<input>
<ID>IN_0</ID>803 </input>
<output>
<ID>OUT_0</ID>629 </output>
<input>
<ID>clock</ID>802 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>61,0.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>814</ID>
<type>AE_SMALL_INVERTER</type>
<position>146.5,-13</position>
<input>
<ID>IN_0</ID>795 </input>
<output>
<ID>OUT_0</ID>804 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>815</ID>
<type>AA_AND2</type>
<position>151.5,-12</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>804 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>61,-1.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>816</ID>
<type>AE_SMALL_INVERTER</type>
<position>165.5,-3.5</position>
<input>
<ID>IN_0</ID>623 </input>
<output>
<ID>OUT_0</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>49</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>69,-2</position>
<output>
<ID>A_greater_B</ID>27 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>107 </input>
<input>
<ID>IN_B_1</ID>108 </input>
<input>
<ID>IN_B_2</ID>109 </input>
<input>
<ID>IN_B_3</ID>110 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_FULLADDER_4BIT</type>
<position>51,21</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>97 </input>
<input>
<ID>IN_B_0</ID>115 </input>
<input>
<ID>IN_B_1</ID>75 </input>
<input>
<ID>IN_B_2</ID>74 </input>
<input>
<ID>IN_B_3</ID>73 </input>
<output>
<ID>OUT_0</ID>111 </output>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>114 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>69,34</position>
<output>
<ID>A_greater_B</ID>28 </output>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_B_0</ID>99 </input>
<input>
<ID>IN_B_1</ID>100 </input>
<input>
<ID>IN_B_2</ID>101 </input>
<input>
<ID>IN_B_3</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>-20,47</position>
<output>
<ID>A_greater_B</ID>1 </output>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>848 </input>
<input>
<ID>IN_2</ID>849 </input>
<input>
<ID>IN_3</ID>850 </input>
<input>
<ID>IN_B_0</ID>843 </input>
<input>
<ID>IN_B_1</ID>844 </input>
<input>
<ID>IN_B_2</ID>845 </input>
<input>
<ID>IN_B_3</ID>846 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_REGISTER4</type>
<position>79,15.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>28 </input>
<input>
<ID>clock</ID>30 </input>
<input>
<ID>load</ID>29 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>78,24.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>CC_PULSE</type>
<position>-70,-18</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>CC_PULSE</type>
<position>78,7.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-73.5,-18</position>
<gparam>LABEL_TEXT pulse</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>78,6</position>
<gparam>LABEL_TEXT update</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>88,16.5</position>
<gparam>LABEL_TEXT blinds</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>-100.5,49</position>
<gparam>LABEL_TEXT outside</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>832</ID>
<type>AA_TOGGLE</type>
<position>-124,87.5</position>
<output>
<ID>OUT_0</ID>853 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>-100,39</position>
<gparam>LABEL_TEXT inside</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>-64,35</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>834</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>-84,83.5</position>
<input>
<ID>ENABLE_0</ID>853 </input>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>852 </input>
<input>
<ID>IN_2</ID>820 </input>
<input>
<ID>IN_3</ID>819 </input>
<output>
<ID>OUT_0</ID>412 </output>
<output>
<ID>OUT_1</ID>409 </output>
<output>
<ID>OUT_2</ID>408 </output>
<output>
<ID>OUT_3</ID>423 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>-57,22</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>-60,35</position>
<input>
<ID>IN_0</ID>850 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>836</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-84,48.5</position>
<input>
<ID>ENABLE_0</ID>853 </input>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>838 </input>
<input>
<ID>IN_2</ID>839 </input>
<input>
<ID>IN_3</ID>840 </input>
<input>
<ID>IN_4</ID>841 </input>
<input>
<ID>IN_5</ID>842 </input>
<input>
<ID>IN_6</ID>836 </input>
<input>
<ID>IN_7</ID>835 </input>
<output>
<ID>OUT_0</ID>850 </output>
<output>
<ID>OUT_1</ID>849 </output>
<output>
<ID>OUT_2</ID>848 </output>
<output>
<ID>OUT_3</ID>847 </output>
<output>
<ID>OUT_4</ID>846 </output>
<output>
<ID>OUT_5</ID>845 </output>
<output>
<ID>OUT_6</ID>844 </output>
<output>
<ID>OUT_7</ID>843 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>-62,29</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>-54,35</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>-50,35</position>
<input>
<ID>IN_0</ID>849 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_OR2</type>
<position>-52,29</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AE_DFF_LOW</type>
<position>-47,22</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>-44,35</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_DFF_LOW</type>
<position>-37,22</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>-40,35</position>
<input>
<ID>IN_0</ID>848 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>844</ID>
<type>AA_LABEL</type>
<position>-95.5,33.5</position>
<gparam>LABEL_TEXT light sensors</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>76</ID>
<type>AE_OR2</type>
<position>-42,29</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>-34,35</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>846</ID>
<type>BA_TRI_STATE</type>
<position>-84.5,115</position>
<input>
<ID>ENABLE_0</ID>853 </input>
<input>
<ID>IN_0</ID>851 </input>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>-27,22</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>-30,35</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>848</ID>
<type>GA_LED</type>
<position>-92,81</position>
<input>
<ID>N_in0</ID>851 </input>
<input>
<ID>N_in1</ID>852 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR2</type>
<position>-32,29</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>849</ID>
<type>AA_LABEL</type>
<position>-134,88.5</position>
<gparam>LABEL_TEXT master</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AE_SMALL_INVERTER</type>
<position>-31,40</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_SMALL_INVERTER</type>
<position>-41,40</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,40</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61,40</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>853</ID>
<type>BA_TRI_STATE</type>
<position>129,33.5</position>
<input>
<ID>ENABLE_0</ID>860 </input>
<input>
<ID>IN_0</ID>854 </input>
<output>
<ID>OUT_0</ID>801 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-80,9</position>
<gparam>LABEL_TEXT shift/load</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>854</ID>
<type>BA_TRI_STATE</type>
<position>129,25</position>
<input>
<ID>ENABLE_0</ID>860 </input>
<input>
<ID>IN_0</ID>855 </input>
<output>
<ID>OUT_0</ID>803 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-75,9</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>855</ID>
<type>AA_LABEL</type>
<position>124.5,118.5</position>
<gparam>LABEL_TEXT sensor</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND2</type>
<position>-64,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>856</ID>
<type>BA_TRI_STATE</type>
<position>129,131</position>
<input>
<ID>ENABLE_0</ID>860 </input>
<input>
<ID>IN_0</ID>859 </input>
<output>
<ID>OUT_0</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_DFF_LOW</type>
<position>-57,-12</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>857</ID>
<type>BA_TRI_STATE</type>
<position>129,125</position>
<input>
<ID>ENABLE_0</ID>860 </input>
<input>
<ID>IN_0</ID>858 </input>
<output>
<ID>OUT_0</ID>433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>-60,1</position>
<input>
<ID>IN_0</ID>846 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AE_OR2</type>
<position>-62,-5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>-54,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>-50,1</position>
<input>
<ID>IN_0</ID>845 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>-52,-5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_DFF_LOW</type>
<position>-47,-12</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND2</type>
<position>-44,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW</type>
<position>-37,-12</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>-40,1</position>
<input>
<ID>IN_0</ID>844 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>-42,-5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND2</type>
<position>-34,1</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_DFF_LOW</type>
<position>-27,-12</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>82 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND2</type>
<position>-30,1</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_OR2</type>
<position>-32,-5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>-31,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>-41,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_SMALL_INVERTER</type>
<position>-61,6</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND2</type>
<position>-14,36</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>-14,30</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>-65,6</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>-65,40</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_SMALL_INVERTER</type>
<position>-19,29</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>-14,20</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>-14,14</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_SMALL_INVERTER</type>
<position>-19,19</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_DFF_LOW</type>
<position>3,31</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_DFF_LOW</type>
<position>11,31</position>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_DFF_LOW</type>
<position>19,31</position>
<input>
<ID>IN_0</ID>74 </input>
<output>
<ID>OUT_0</ID>75 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_DFF_LOW</type>
<position>27,31</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>115 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>-5,33</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_DFF_LOW</type>
<position>3,15</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>77 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_DFF_LOW</type>
<position>11.5,15</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>78 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_DFF_LOW</type>
<position>19.5,15</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_DFF_LOW</type>
<position>27.5,15</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_OR2</type>
<position>-5,17</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>-29,128.5</position>
<gparam>LABEL_TEXT loop activate-able</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>-91.5,115</position>
<output>
<ID>OUT_0</ID>851 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-6,110.5</position>
<gparam>LABEL_TEXT device 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-6,97.5</position>
<gparam>LABEL_TEXT device 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_REGISTER4</type>
<position>-59,104</position>
<output>
<ID>OUT_0</ID>121 </output>
<output>
<ID>OUT_1</ID>120 </output>
<output>
<ID>OUT_2</ID>119 </output>
<output>
<ID>OUT_3</ID>118 </output>
<input>
<ID>clear</ID>131 </input>
<input>
<ID>clock</ID>123 </input>
<input>
<ID>count_enable</ID>125 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND4</type>
<position>-50,104.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>121 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>131</ID>
<type>BE_NOR2</type>
<position>-14,115.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>BB_CLOCK</type>
<position>-66,98</position>
<output>
<ID>CLK</ID>123 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 1</lparam></gate>
<gate>
<ID>133</ID>
<type>BE_NOR2</type>
<position>-14,108.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>-8,108.5</position>
<input>
<ID>N_in0</ID>116 </input>
<input>
<ID>N_in1</ID>860 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>BE_NOR2</type>
<position>-68,111</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>BE_NOR2</type>
<position>-68,104</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>BE_NOR2</type>
<position>-40,108</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>BE_NOR2</type>
<position>-40,101</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AE_SMALL_INVERTER</type>
<position>-75,103</position>
<input>
<ID>IN_0</ID>139 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>-97,115</position>
<gparam>LABEL_TEXT occ. sensor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>-29,126</position>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_OR2</type>
<position>-74,112</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_OR2</type>
<position>-58,95</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>-22,114</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>-22,110</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>-14,102.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>BE_NOR2</type>
<position>-14,95.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>-8,95.5</position>
<input>
<ID>N_in0</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>-22,101</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>-22,97</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_SMALL_INVERTER</type>
<position>-27,120</position>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_TOGGLE</type>
<position>-92,85</position>
<output>
<ID>OUT_0</ID>819 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_TOGGLE</type>
<position>-92,83</position>
<output>
<ID>OUT_0</ID>820 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>407</ID>
<type>AE_OR2</type>
<position>-67,79</position>
<input>
<ID>IN_0</ID>408 </input>
<input>
<ID>IN_1</ID>409 </input>
<output>
<ID>OUT</ID>410 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>-59,78</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>413 </input>
<output>
<ID>OUT</ID>411 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_TOGGLE</type>
<position>-92,79</position>
<output>
<ID>OUT_0</ID>822 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>410</ID>
<type>AE_OR2</type>
<position>-51,84</position>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>411 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>AA_LABEL</type>
<position>-97,85</position>
<gparam>LABEL_TEXT mag. lock</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>412</ID>
<type>AA_LABEL</type>
<position>-98.5,83</position>
<gparam>LABEL_TEXT sound sensor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AA_LABEL</type>
<position>-95,79</position>
<gparam>LABEL_TEXT GPS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>AA_INVERTER</type>
<position>-67,71</position>
<input>
<ID>IN_0</ID>412 </input>
<output>
<ID>OUT_0</ID>413 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>416</ID>
<type>BE_NOR2</type>
<position>-43,83</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>418 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>BE_NOR2</type>
<position>-43,76</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>-77.5,62</position>
<gparam>LABEL_TEXT reset</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>CC_PULSE</type>
<position>-74,62</position>
<output>
<ID>OUT_0</ID>417 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>GA_LED</type>
<position>-34,76</position>
<input>
<ID>N_in0</ID>418 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>421</ID>
<type>AA_LABEL</type>
<position>-22.5,76</position>
<gparam>LABEL_TEXT alarm, police, video, notify</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>GA_LED</type>
<position>-20,61</position>
<input>
<ID>N_in0</ID>422 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>BE_NOR2</type>
<position>-27,68</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>422 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>424</ID>
<type>BE_NOR2</type>
<position>-27,61</position>
<input>
<ID>IN_0</ID>424 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>422 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>CC_PULSE</type>
<position>-50,64</position>
<output>
<ID>OUT_0</ID>416 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AE_OR2</type>
<position>-43,63</position>
<input>
<ID>IN_0</ID>416 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>421 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>427</ID>
<type>AA_LABEL</type>
<position>-54.5,64</position>
<gparam>LABEL_TEXT hang up</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_LABEL</type>
<position>-14,61</position>
<gparam>LABEL_TEXT conversation</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_AND2</type>
<position>-35,69</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>CC_PULSE</type>
<position>-50,68</position>
<output>
<ID>OUT_0</ID>419 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_LABEL</type>
<position>-52.5,68</position>
<gparam>LABEL_TEXT call</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>432</ID>
<type>AA_TOGGLE</type>
<position>177.5,108</position>
<output>
<ID>OUT_0</ID>489 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>433</ID>
<type>AA_LABEL</type>
<position>177.5,106.5</position>
<gparam>LABEL_TEXT Reset</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>164,153</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>168.5,116.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AA_TOGGLE</type>
<position>123,131</position>
<output>
<ID>OUT_0</ID>859 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>124,121</position>
<gparam>LABEL_TEXT temperature</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>162,107.5</position>
<gparam>LABEL_TEXT Update</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>114.5,131.5</position>
<gparam>LABEL_TEXT Increase/Decrease</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>AE_SMALL_INVERTER</type>
<position>176.5,124</position>
<input>
<ID>IN_0</ID>433 </input>
<output>
<ID>OUT_0</ID>434 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_LABEL</type>
<position>119,125</position>
<gparam>LABEL_TEXT On/Off</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>443</ID>
<type>AA_TOGGLE</type>
<position>123,125</position>
<output>
<ID>OUT_0</ID>858 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>444</ID>
<type>AE_REGISTER8</type>
<position>176.5,116</position>
<output>
<ID>OUT_0</ID>443 </output>
<output>
<ID>OUT_1</ID>442 </output>
<output>
<ID>OUT_2</ID>441 </output>
<output>
<ID>OUT_3</ID>440 </output>
<output>
<ID>OUT_4</ID>439 </output>
<output>
<ID>OUT_5</ID>438 </output>
<output>
<ID>OUT_6</ID>437 </output>
<output>
<ID>OUT_7</ID>436 </output>
<output>
<ID>carry_out</ID>477 </output>
<input>
<ID>clear</ID>489 </input>
<input>
<ID>clock</ID>857 </input>
<input>
<ID>count_enable</ID>434 </input>
<input>
<ID>count_up</ID>435 </input>
<input>
<ID>load</ID>433 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_LABEL</type>
<position>189,187.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>446</ID>
<type>BB_CLOCK</type>
<position>167.5,107.5</position>
<output>
<ID>CLK</ID>857 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>447</ID>
<type>BE_JKFF_LOW</type>
<position>145.5,143</position>
<input>
<ID>J</ID>476 </input>
<input>
<ID>K</ID>476 </input>
<output>
<ID>Q</ID>533 </output>
<input>
<ID>clock</ID>477 </input>
<output>
<ID>nQ</ID>480 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>448</ID>
<type>BE_JKFF_LOW</type>
<position>170.5,143</position>
<input>
<ID>J</ID>484 </input>
<input>
<ID>K</ID>484 </input>
<output>
<ID>Q</ID>517 </output>
<input>
<ID>clock</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>449</ID>
<type>AA_TOGGLE</type>
<position>136.5,143</position>
<output>
<ID>OUT_0</ID>476 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_LABEL</type>
<position>133,143</position>
<gparam>LABEL_TEXT logic1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>451</ID>
<type>AA_AND2</type>
<position>153.5,148</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>533 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>AA_AND2</type>
<position>153.5,138</position>
<input>
<ID>IN_0</ID>480 </input>
<input>
<ID>IN_1</ID>478 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>453</ID>
<type>AE_SMALL_INVERTER</type>
<position>146.5,137</position>
<input>
<ID>IN_0</ID>435 </input>
<output>
<ID>OUT_0</ID>478 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>454</ID>
<type>AE_OR2</type>
<position>161.5,143</position>
<input>
<ID>IN_0</ID>482 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>484 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>239,166</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>262,115.5</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_LABEL</type>
<position>239,64.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>AE_OR2</type>
<position>240.5,129</position>
<input>
<ID>IN_0</ID>474 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>455 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>459</ID>
<type>AE_OR2</type>
<position>240.5,125</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>472 </input>
<output>
<ID>OUT</ID>454 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AE_OR2</type>
<position>240.5,121</position>
<input>
<ID>IN_0</ID>479 </input>
<input>
<ID>IN_1</ID>471 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_OR2</type>
<position>240.5,117</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>470 </input>
<output>
<ID>OUT</ID>452 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>AE_OR2</type>
<position>240.5,113</position>
<input>
<ID>IN_0</ID>485 </input>
<input>
<ID>IN_1</ID>469 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>AE_OR2</type>
<position>240.5,109</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>468 </input>
<output>
<ID>OUT</ID>450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>AE_OR2</type>
<position>240.5,105</position>
<input>
<ID>IN_0</ID>487 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>449 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>465</ID>
<type>AE_OR2</type>
<position>240.5,101</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>466 </input>
<output>
<ID>OUT</ID>448 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>466</ID>
<type>AA_AND2</type>
<position>217.5,180</position>
<input>
<ID>IN_0</ID>491 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>465 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>467</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,181</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>491 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND2</type>
<position>217.5,176</position>
<input>
<ID>IN_0</ID>506 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND2</type>
<position>217.5,172</position>
<input>
<ID>IN_0</ID>505 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>463 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_AND2</type>
<position>217.5,168</position>
<input>
<ID>IN_0</ID>504 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_AND2</type>
<position>217.5,164</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>496 </input>
<output>
<ID>OUT</ID>461 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_AND2</type>
<position>217.5,160</position>
<input>
<ID>IN_0</ID>502 </input>
<input>
<ID>IN_1</ID>497 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>AA_AND2</type>
<position>217.5,156</position>
<input>
<ID>IN_0</ID>501 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>459 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>474</ID>
<type>AA_AND2</type>
<position>217.5,152</position>
<input>
<ID>IN_0</ID>500 </input>
<input>
<ID>IN_1</ID>499 </input>
<output>
<ID>OUT</ID>458 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_AND2</type>
<position>217.5,146</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>492 </input>
<output>
<ID>OUT</ID>474 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>AA_AND2</type>
<position>217.5,142</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>493 </input>
<output>
<ID>OUT</ID>475 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>477</ID>
<type>AA_AND2</type>
<position>217.5,138</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>AA_AND2</type>
<position>217.5,134</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>481 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>479</ID>
<type>AA_AND2</type>
<position>217.5,130</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>496 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>217.5,126</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>497 </input>
<output>
<ID>OUT</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>AA_AND2</type>
<position>217.5,122</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>482</ID>
<type>AA_AND2</type>
<position>217.5,118</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>499 </input>
<output>
<ID>OUT</ID>488 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>483</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,177</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>484</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,173</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>485</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,169</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>486</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,165</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>503 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>487</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,161</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>488</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,157</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>501 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>489</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,153</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>500 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_AND2</type>
<position>217.5,112</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>508 </input>
<output>
<ID>OUT</ID>473 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>491</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,113</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_AND2</type>
<position>217.5,108</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>509 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_AND2</type>
<position>217.5,104</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>217.5,100</position>
<input>
<ID>IN_0</ID>521 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>470 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_AND2</type>
<position>217.5,96</position>
<input>
<ID>IN_0</ID>520 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>469 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>496</ID>
<type>AA_AND2</type>
<position>217.5,92</position>
<input>
<ID>IN_0</ID>519 </input>
<input>
<ID>IN_1</ID>513 </input>
<output>
<ID>OUT</ID>468 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>497</ID>
<type>AA_AND2</type>
<position>217.5,88</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>514 </input>
<output>
<ID>OUT</ID>467 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>498</ID>
<type>AA_AND2</type>
<position>217.5,84</position>
<input>
<ID>IN_0</ID>516 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_AND2</type>
<position>217.5,78</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>508 </input>
<output>
<ID>OUT</ID>445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>AA_AND2</type>
<position>217.5,74</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>509 </input>
<output>
<ID>OUT</ID>444 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_AND2</type>
<position>217.5,70</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>510 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>502</ID>
<type>AA_AND2</type>
<position>217.5,66</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>511 </input>
<output>
<ID>OUT</ID>431 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_AND2</type>
<position>217.5,62</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AA_AND2</type>
<position>217.5,58</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>513 </input>
<output>
<ID>OUT</ID>429 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>505</ID>
<type>AA_AND2</type>
<position>217.5,54</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>514 </input>
<output>
<ID>OUT</ID>428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_AND2</type>
<position>217.5,50</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>515 </input>
<output>
<ID>OUT</ID>427 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>507</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,109</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>508</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,105</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>509</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,101</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>510</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,97</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>511</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,93</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>519 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>512</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,89</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>513</ID>
<type>AE_SMALL_INVERTER</type>
<position>212.5,85</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_LABEL</type>
<position>196,183</position>
<gparam>LABEL_TEXT ~D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>515</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,178</position>
<input>
<ID>IN_0</ID>443 </input>
<output>
<ID>OUT_0</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>516</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,174</position>
<input>
<ID>IN_0</ID>442 </input>
<output>
<ID>OUT_0</ID>525 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>517</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,170</position>
<input>
<ID>IN_0</ID>441 </input>
<output>
<ID>OUT_0</ID>526 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>518</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,166</position>
<input>
<ID>IN_0</ID>440 </input>
<output>
<ID>OUT_0</ID>527 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>519</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,162</position>
<input>
<ID>IN_0</ID>439 </input>
<output>
<ID>OUT_0</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>520</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,158</position>
<input>
<ID>IN_0</ID>438 </input>
<output>
<ID>OUT_0</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>521</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,154</position>
<input>
<ID>IN_0</ID>437 </input>
<output>
<ID>OUT_0</ID>530 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>522</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,150</position>
<input>
<ID>IN_0</ID>436 </input>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>523</ID>
<type>AE_OR2</type>
<position>197.5,179</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>524 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>524</ID>
<type>AE_OR2</type>
<position>197.5,175</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>525 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>525</ID>
<type>AE_OR2</type>
<position>197.5,171</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>526 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>526</ID>
<type>AE_OR2</type>
<position>197.5,167</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>527 </input>
<output>
<ID>OUT</ID>495 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>AE_OR2</type>
<position>197.5,163</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>528 </input>
<output>
<ID>OUT</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>AE_OR2</type>
<position>197.5,159</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>529 </input>
<output>
<ID>OUT</ID>497 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>529</ID>
<type>AE_OR2</type>
<position>197.5,155</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>530 </input>
<output>
<ID>OUT</ID>498 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>530</ID>
<type>AE_OR2</type>
<position>197.5,151</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>531 </input>
<output>
<ID>OUT</ID>499 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>531</ID>
<type>AE_SMALL_INVERTER</type>
<position>178.5,180</position>
<input>
<ID>IN_0</ID>533 </input>
<output>
<ID>OUT_0</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>532</ID>
<type>AA_LABEL</type>
<position>197,115</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>533</ID>
<type>AE_OR2</type>
<position>197.5,111</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>443 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>534</ID>
<type>AE_OR2</type>
<position>197.5,107</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>535</ID>
<type>AE_OR2</type>
<position>197.5,103</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>441 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>536</ID>
<type>AE_OR2</type>
<position>197.5,99</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>440 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AE_OR2</type>
<position>197.5,95</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>439 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>538</ID>
<type>AE_OR2</type>
<position>197.5,91</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>438 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>AE_OR2</type>
<position>197.5,87</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>437 </input>
<output>
<ID>OUT</ID>514 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>540</ID>
<type>AE_OR2</type>
<position>197.5,83</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>515 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>541</ID>
<type>AE_REGISTER8</type>
<position>233.5,165.5</position>
<input>
<ID>IN_0</ID>465 </input>
<input>
<ID>IN_1</ID>464 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>462 </input>
<input>
<ID>IN_4</ID>461 </input>
<input>
<ID>IN_5</ID>460 </input>
<input>
<ID>IN_6</ID>459 </input>
<input>
<ID>IN_7</ID>458 </input>
<input>
<ID>clock</ID>457 </input>
<input>
<ID>load</ID>456 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>542</ID>
<type>AE_REGISTER8</type>
<position>233.5,63.5</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>444 </input>
<input>
<ID>IN_2</ID>432 </input>
<input>
<ID>IN_3</ID>431 </input>
<input>
<ID>IN_4</ID>430 </input>
<input>
<ID>IN_5</ID>429 </input>
<input>
<ID>IN_6</ID>428 </input>
<input>
<ID>IN_7</ID>427 </input>
<input>
<ID>clock</ID>425 </input>
<input>
<ID>load</ID>426 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>543</ID>
<type>BB_CLOCK</type>
<position>232.5,54.5</position>
<output>
<ID>CLK</ID>425 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>544</ID>
<type>BB_CLOCK</type>
<position>232.5,156.5</position>
<output>
<ID>CLK</ID>457 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>545</ID>
<type>AA_TOGGLE</type>
<position>232.5,173.5</position>
<output>
<ID>OUT_0</ID>456 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>546</ID>
<type>AE_REGISTER8</type>
<position>256.5,114.5</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>454 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>452 </input>
<input>
<ID>IN_4</ID>451 </input>
<input>
<ID>IN_5</ID>450 </input>
<input>
<ID>IN_6</ID>449 </input>
<input>
<ID>IN_7</ID>448 </input>
<input>
<ID>clock</ID>447 </input>
<input>
<ID>load</ID>446 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>547</ID>
<type>BB_CLOCK</type>
<position>255.5,105.5</position>
<output>
<ID>CLK</ID>447 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>548</ID>
<type>AA_TOGGLE</type>
<position>255.5,122.5</position>
<output>
<ID>OUT_0</ID>446 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>549</ID>
<type>AA_TOGGLE</type>
<position>232.5,71.5</position>
<output>
<ID>OUT_0</ID>426 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>550</ID>
<type>AA_AND2</type>
<position>156,-19</position>
<input>
<ID>IN_0</ID>590 </input>
<input>
<ID>IN_1</ID>622 </input>
<output>
<ID>OUT</ID>589 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>551</ID>
<type>AA_TOGGLE</type>
<position>123,25</position>
<output>
<ID>OUT_0</ID>855 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>552</ID>
<type>AE_SMALL_INVERTER</type>
<position>337,-9.5</position>
<input>
<ID>IN_0</ID>799 </input>
<output>
<ID>OUT_0</ID>805 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>553</ID>
<type>AA_LABEL</type>
<position>116.5,25</position>
<gparam>LABEL_TEXT Change Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>554</ID>
<type>AE_SMALL_INVERTER</type>
<position>339,-92.5</position>
<input>
<ID>IN_0</ID>800 </input>
<output>
<ID>OUT_0</ID>806 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>556</ID>
<type>AA_AND4</type>
<position>281.5,24</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>714 </input>
<output>
<ID>OUT</ID>811 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND4</type>
<position>281.5,16</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>796 </input>
<output>
<ID>OUT</ID>812 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_AND4</type>
<position>281.5,8</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>562</ID>
<type>AA_AND4</type>
<position>281.5,0</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>564</ID>
<type>AA_AND4</type>
<position>281.5,-8</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>566</ID>
<type>AA_AND4</type>
<position>281.5,-16</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>568</ID>
<type>AA_AND4</type>
<position>281.5,-24</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>570</ID>
<type>AA_AND4</type>
<position>281.5,-32</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_AND2</type>
<position>170,-37</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>626 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>AE_SMALL_INVERTER</type>
<position>273.5,35</position>
<input>
<ID>IN_0</ID>798 </input>
<output>
<ID>OUT_0</ID>740 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>574</ID>
<type>AE_SMALL_INVERTER</type>
<position>275.5,35</position>
<input>
<ID>IN_0</ID>797 </input>
<output>
<ID>OUT_0</ID>719 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>575</ID>
<type>AA_AND4</type>
<position>281.5,-50.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>714 </input>
<output>
<ID>OUT</ID>799 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>576</ID>
<type>AE_SMALL_INVERTER</type>
<position>277.5,35</position>
<input>
<ID>IN_0</ID>796 </input>
<output>
<ID>OUT_0</ID>714 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>577</ID>
<type>AE_DFF_LOW</type>
<position>181.5,-13</position>
<input>
<ID>IN_0</ID>566 </input>
<output>
<ID>OUT_0</ID>547 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>578</ID>
<type>AA_AND2</type>
<position>184,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>543 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>579</ID>
<type>AE_SMALL_INVERTER</type>
<position>141,-22</position>
<input>
<ID>IN_0</ID>795 </input>
<output>
<ID>OUT_0</ID>660 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>580</ID>
<type>AA_AND2</type>
<position>188,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>567 </input>
<output>
<ID>OUT</ID>544 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>581</ID>
<type>AE_OR2</type>
<position>186,-6</position>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>543 </input>
<output>
<ID>OUT</ID>568 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>582</ID>
<type>AE_SMALL_INVERTER</type>
<position>141,-26</position>
<input>
<ID>IN_0</ID>660 </input>
<output>
<ID>OUT_0</ID>585 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>583</ID>
<type>AE_OR2</type>
<position>163.5,-30.5</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>586 </input>
<output>
<ID>OUT</ID>587 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>584</ID>
<type>AE_SMALL_INVERTER</type>
<position>178.5,3.5</position>
<input>
<ID>IN_0</ID>700 </input>
<output>
<ID>OUT_0</ID>661 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>585</ID>
<type>AE_DFF_LOW</type>
<position>190.5,-13</position>
<input>
<ID>IN_0</ID>568 </input>
<output>
<ID>OUT_0</ID>550 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>586</ID>
<type>AE_SMALL_INVERTER</type>
<position>155.5,-40</position>
<input>
<ID>IN_0</ID>585 </input>
<output>
<ID>OUT_0</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>587</ID>
<type>AA_AND2</type>
<position>193,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>550 </input>
<output>
<ID>OUT</ID>548 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>588</ID>
<type>AA_AND2</type>
<position>197,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>580 </input>
<output>
<ID>OUT</ID>549 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>589</ID>
<type>AE_OR2</type>
<position>195,-6</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>548 </input>
<output>
<ID>OUT</ID>570 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>590</ID>
<type>AE_DFF_LOW</type>
<position>199.5,-13</position>
<input>
<ID>IN_0</ID>570 </input>
<output>
<ID>OUT_0</ID>553 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>591</ID>
<type>AA_AND2</type>
<position>202,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>553 </input>
<output>
<ID>OUT</ID>551 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>592</ID>
<type>AA_AND2</type>
<position>206,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>579 </input>
<output>
<ID>OUT</ID>552 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>593</ID>
<type>AE_OR2</type>
<position>204,-6</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>551 </input>
<output>
<ID>OUT</ID>569 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>594</ID>
<type>AE_DFF_LOW</type>
<position>209,-13</position>
<input>
<ID>IN_0</ID>569 </input>
<output>
<ID>OUT_0</ID>556 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>595</ID>
<type>AA_AND2</type>
<position>211.5,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>556 </input>
<output>
<ID>OUT</ID>554 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>596</ID>
<type>AA_AND2</type>
<position>215.5,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>578 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AE_OR2</type>
<position>213.5,-6</position>
<input>
<ID>IN_0</ID>555 </input>
<input>
<ID>IN_1</ID>554 </input>
<output>
<ID>OUT</ID>571 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>598</ID>
<type>AE_DFF_LOW</type>
<position>218,-13</position>
<input>
<ID>IN_0</ID>571 </input>
<output>
<ID>OUT_0</ID>559 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_AND2</type>
<position>220.5,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>559 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_AND2</type>
<position>224.5,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>577 </input>
<output>
<ID>OUT</ID>558 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AE_OR2</type>
<position>222.5,-6</position>
<input>
<ID>IN_0</ID>558 </input>
<input>
<ID>IN_1</ID>557 </input>
<output>
<ID>OUT</ID>572 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>AE_DFF_LOW</type>
<position>227,-13</position>
<input>
<ID>IN_0</ID>572 </input>
<output>
<ID>OUT_0</ID>562 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_AND2</type>
<position>229.5,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>562 </input>
<output>
<ID>OUT</ID>560 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>604</ID>
<type>AA_AND2</type>
<position>233.5,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>576 </input>
<output>
<ID>OUT</ID>561 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>605</ID>
<type>AE_OR2</type>
<position>231.5,-6</position>
<input>
<ID>IN_0</ID>561 </input>
<input>
<ID>IN_1</ID>560 </input>
<output>
<ID>OUT</ID>573 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>606</ID>
<type>AE_DFF_LOW</type>
<position>236,-13</position>
<input>
<ID>IN_0</ID>573 </input>
<output>
<ID>OUT_0</ID>565 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_AND2</type>
<position>238.5,0</position>
<input>
<ID>IN_0</ID>663 </input>
<input>
<ID>IN_1</ID>565 </input>
<output>
<ID>OUT</ID>563 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_AND2</type>
<position>242.5,0</position>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>575 </input>
<output>
<ID>OUT</ID>564 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>609</ID>
<type>AE_OR2</type>
<position>240.5,-6</position>
<input>
<ID>IN_0</ID>564 </input>
<input>
<ID>IN_1</ID>563 </input>
<output>
<ID>OUT</ID>574 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>611</ID>
<type>AE_DFF_LOW</type>
<position>245,-13</position>
<input>
<ID>IN_0</ID>574 </input>
<output>
<ID>OUT_0</ID>542 </output>
<input>
<ID>clock</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>612</ID>
<type>AA_AND4</type>
<position>281.5,-58.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>796 </input>
<output>
<ID>OUT</ID>800 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>613</ID>
<type>AE_REGISTER8</type>
<position>168.5,9.5</position>
<input>
<ID>IN_0</ID>619 </input>
<input>
<ID>IN_1</ID>620 </input>
<input>
<ID>IN_2</ID>618 </input>
<input>
<ID>IN_3</ID>617 </input>
<input>
<ID>IN_4</ID>616 </input>
<input>
<ID>IN_5</ID>615 </input>
<input>
<ID>IN_6</ID>614 </input>
<input>
<ID>IN_7</ID>613 </input>
<output>
<ID>OUT_0</ID>566 </output>
<output>
<ID>OUT_1</ID>567 </output>
<output>
<ID>OUT_2</ID>580 </output>
<output>
<ID>OUT_3</ID>579 </output>
<output>
<ID>OUT_4</ID>578 </output>
<output>
<ID>OUT_5</ID>577 </output>
<output>
<ID>OUT_6</ID>576 </output>
<output>
<ID>OUT_7</ID>575 </output>
<input>
<ID>clock</ID>665 </input>
<input>
<ID>load</ID>621 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>615</ID>
<type>BB_CLOCK</type>
<position>151,-37</position>
<output>
<ID>CLK</ID>582 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_AND2</type>
<position>158,-34.5</position>
<input>
<ID>IN_0</ID>584 </input>
<input>
<ID>IN_1</ID>582 </input>
<output>
<ID>OUT</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_REGISTER4</type>
<position>156.5,-26.5</position>
<output>
<ID>OUT_0</ID>622 </output>
<output>
<ID>OUT_3</ID>590 </output>
<input>
<ID>clear</ID>589 </input>
<input>
<ID>clock</ID>587 </input>
<input>
<ID>count_enable</ID>588 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>618</ID>
<type>AA_TOGGLE</type>
<position>149.5,-26.5</position>
<output>
<ID>OUT_0</ID>588 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>619</ID>
<type>AE_SMALL_INVERTER</type>
<position>146.5,-31.5</position>
<input>
<ID>IN_0</ID>589 </input>
<output>
<ID>OUT_0</ID>583 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>620</ID>
<type>AA_AND2</type>
<position>151.5,-32.5</position>
<input>
<ID>IN_0</ID>583 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>621</ID>
<type>AE_REGISTER8</type>
<position>338,-2.5</position>
<input>
<ID>IN_0</ID>592 </input>
<input>
<ID>IN_1</ID>593 </input>
<input>
<ID>IN_2</ID>594 </input>
<input>
<ID>IN_3</ID>595 </input>
<input>
<ID>IN_4</ID>596 </input>
<input>
<ID>IN_5</ID>597 </input>
<input>
<ID>IN_6</ID>598 </input>
<input>
<ID>IN_7</ID>599 </input>
<output>
<ID>OUT_0</ID>777 </output>
<output>
<ID>OUT_1</ID>778 </output>
<output>
<ID>OUT_2</ID>779 </output>
<output>
<ID>OUT_3</ID>780 </output>
<output>
<ID>OUT_4</ID>781 </output>
<output>
<ID>OUT_5</ID>807 </output>
<output>
<ID>OUT_6</ID>783 </output>
<output>
<ID>OUT_7</ID>784 </output>
<input>
<ID>clock</ID>805 </input>
<input>
<ID>load</ID>601 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 210</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>622</ID>
<type>AE_DFF_LOW</type>
<position>311,-28.5</position>
<input>
<ID>IN_0</ID>811 </input>
<output>
<ID>OUT_0</ID>592 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>623</ID>
<type>AE_DFF_LOW</type>
<position>311,-20</position>
<input>
<ID>IN_0</ID>592 </input>
<output>
<ID>OUT_0</ID>593 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>624</ID>
<type>AE_DFF_LOW</type>
<position>311,-11.5</position>
<input>
<ID>IN_0</ID>593 </input>
<output>
<ID>OUT_0</ID>594 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>625</ID>
<type>AE_DFF_LOW</type>
<position>311,-3.5</position>
<input>
<ID>IN_0</ID>594 </input>
<output>
<ID>OUT_0</ID>595 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>626</ID>
<type>AE_DFF_LOW</type>
<position>311,4</position>
<input>
<ID>IN_0</ID>595 </input>
<output>
<ID>OUT_0</ID>596 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>627</ID>
<type>AE_DFF_LOW</type>
<position>311,11.5</position>
<input>
<ID>IN_0</ID>596 </input>
<output>
<ID>OUT_0</ID>597 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>628</ID>
<type>AE_DFF_LOW</type>
<position>311,19</position>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>598 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>629</ID>
<type>AE_DFF_LOW</type>
<position>311,26.5</position>
<input>
<ID>IN_0</ID>598 </input>
<output>
<ID>OUT_0</ID>599 </output>
<input>
<ID>clock</ID>799 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>630</ID>
<type>AA_AND4</type>
<position>281.5,-66.5</position>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>631</ID>
<type>AA_TOGGLE</type>
<position>337,5.5</position>
<output>
<ID>OUT_0</ID>601 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>632</ID>
<type>AE_REGISTER8</type>
<position>340,-85.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>604 </input>
<input>
<ID>IN_2</ID>605 </input>
<input>
<ID>IN_3</ID>606 </input>
<input>
<ID>IN_4</ID>607 </input>
<input>
<ID>IN_5</ID>608 </input>
<input>
<ID>IN_6</ID>609 </input>
<input>
<ID>IN_7</ID>610 </input>
<output>
<ID>OUT_0</ID>785 </output>
<output>
<ID>OUT_1</ID>786 </output>
<output>
<ID>OUT_2</ID>787 </output>
<output>
<ID>OUT_3</ID>788 </output>
<output>
<ID>OUT_4</ID>789 </output>
<output>
<ID>OUT_5</ID>790 </output>
<output>
<ID>OUT_6</ID>791 </output>
<output>
<ID>OUT_7</ID>776 </output>
<input>
<ID>clock</ID>806 </input>
<input>
<ID>load</ID>612 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 18</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>633</ID>
<type>AE_DFF_LOW</type>
<position>313,-111.5</position>
<input>
<ID>IN_0</ID>812 </input>
<output>
<ID>OUT_0</ID>603 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>634</ID>
<type>AE_DFF_LOW</type>
<position>313,-103</position>
<input>
<ID>IN_0</ID>603 </input>
<output>
<ID>OUT_0</ID>604 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>635</ID>
<type>AE_DFF_LOW</type>
<position>313,-95</position>
<input>
<ID>IN_0</ID>604 </input>
<output>
<ID>OUT_0</ID>605 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>636</ID>
<type>AE_DFF_LOW</type>
<position>313,-87</position>
<input>
<ID>IN_0</ID>605 </input>
<output>
<ID>OUT_0</ID>606 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>637</ID>
<type>AE_DFF_LOW</type>
<position>313,-79</position>
<input>
<ID>IN_0</ID>606 </input>
<output>
<ID>OUT_0</ID>607 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>638</ID>
<type>AE_DFF_LOW</type>
<position>313,-71</position>
<input>
<ID>IN_0</ID>607 </input>
<output>
<ID>OUT_0</ID>608 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>639</ID>
<type>AE_DFF_LOW</type>
<position>313,-63</position>
<input>
<ID>IN_0</ID>608 </input>
<output>
<ID>OUT_0</ID>609 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>640</ID>
<type>AE_DFF_LOW</type>
<position>313,-55</position>
<input>
<ID>IN_0</ID>609 </input>
<output>
<ID>OUT_0</ID>610 </output>
<input>
<ID>clock</ID>800 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>641</ID>
<type>AA_AND2</type>
<position>160.5,-11</position>
<input>
<ID>IN_0</ID>629 </input>
<input>
<ID>IN_1</ID>611 </input>
<output>
<ID>OUT</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>642</ID>
<type>AA_TOGGLE</type>
<position>339,-77.5</position>
<output>
<ID>OUT_0</ID>612 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>643</ID>
<type>AA_TOGGLE</type>
<position>141.5,15.5</position>
<output>
<ID>OUT_0</ID>613 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>644</ID>
<type>AA_TOGGLE</type>
<position>141.5,13.5</position>
<output>
<ID>OUT_0</ID>614 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>645</ID>
<type>AA_TOGGLE</type>
<position>141.5,11.5</position>
<output>
<ID>OUT_0</ID>615 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>646</ID>
<type>AA_TOGGLE</type>
<position>141.5,9.5</position>
<output>
<ID>OUT_0</ID>616 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>647</ID>
<type>AA_TOGGLE</type>
<position>141.5,7.5</position>
<output>
<ID>OUT_0</ID>617 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>648</ID>
<type>AA_TOGGLE</type>
<position>141.5,5.5</position>
<output>
<ID>OUT_0</ID>618 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_TOGGLE</type>
<position>141.5,3.5</position>
<output>
<ID>OUT_0</ID>620 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>650</ID>
<type>AA_TOGGLE</type>
<position>141.5,1.5</position>
<output>
<ID>OUT_0</ID>619 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>651</ID>
<type>AA_TOGGLE</type>
<position>167.5,17.5</position>
<output>
<ID>OUT_0</ID>621 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_LABEL</type>
<position>135.5,8.5</position>
<gparam>LABEL_TEXT New Color</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>653</ID>
<type>AA_AND2</type>
<position>178,-36</position>
<input>
<ID>IN_0</ID>629 </input>
<input>
<ID>IN_1</ID>626 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>655</ID>
<type>AE_OR2</type>
<position>149,-4.5</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>629 </input>
<output>
<ID>OUT</ID>795 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>AA_AND2</type>
<position>178,-44.5</position>
<input>
<ID>IN_0</ID>626 </input>
<input>
<ID>IN_1</ID>810 </input>
<output>
<ID>OUT</ID>581 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_AND2</type>
<position>187.5,-30.5</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>611 </input>
<output>
<ID>OUT</ID>662 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>AA_AND4</type>
<position>281.5,-74.5</position>
<input>
<ID>IN_1</ID>740 </input>
<input>
<ID>IN_2</ID>797 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>659</ID>
<type>AE_SMALL_INVERTER</type>
<position>204,-27</position>
<input>
<ID>IN_0</ID>658 </input>
<output>
<ID>OUT_0</ID>546 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>660</ID>
<type>AI_MUX_8x1</type>
<position>453.5,-57.5</position>
<input>
<ID>IN_0</ID>809 </input>
<input>
<ID>IN_1</ID>808 </input>
<output>
<ID>OUT</ID>625 </output>
<input>
<ID>SEL_0</ID>796 </input>
<input>
<ID>SEL_1</ID>797 </input>
<input>
<ID>SEL_2</ID>798 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>661</ID>
<type>AA_MUX_2x1</type>
<position>562.5,-71.5</position>
<input>
<ID>IN_0</ID>774 </input>
<input>
<ID>IN_1</ID>625 </input>
<output>
<ID>OUT</ID>764 </output>
<input>
<ID>SEL_0</ID>810 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_LABEL</type>
<position>566,-85</position>
<gparam>LABEL_TEXT Default lights</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>663</ID>
<type>AA_LABEL</type>
<position>533.5,-69</position>
<gparam>LABEL_TEXT Notification lights</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>664</ID>
<type>AA_LABEL</type>
<position>596,-37.5</position>
<gparam>LABEL_TEXT Light</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>665</ID>
<type>AE_DFF_LOW</type>
<position>377,-85</position>
<input>
<ID>IN_0</ID>785 </input>
<output>
<ID>OUT_0</ID>630 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>666</ID>
<type>AA_AND2</type>
<position>379.5,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>630 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_AND2</type>
<position>383.5,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>786 </input>
<output>
<ID>OUT</ID>628 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>668</ID>
<type>AE_OR2</type>
<position>381.5,-78</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>627 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>669</ID>
<type>AA_AND2</type>
<position>205,-30.5</position>
<input>
<ID>IN_0</ID>658 </input>
<input>
<ID>IN_1</ID>658 </input>
<output>
<ID>OUT</ID>782 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>AE_SMALL_INVERTER</type>
<position>198.5,-30.5</position>
<input>
<ID>IN_0</ID>662 </input>
<output>
<ID>OUT_0</ID>658 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>671</ID>
<type>AE_DFF_LOW</type>
<position>386,-85</position>
<input>
<ID>IN_0</ID>651 </input>
<output>
<ID>OUT_0</ID>633 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>672</ID>
<type>AA_AND2</type>
<position>388.5,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>633 </input>
<output>
<ID>OUT</ID>631 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>673</ID>
<type>AA_AND2</type>
<position>392.5,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>787 </input>
<output>
<ID>OUT</ID>632 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>674</ID>
<type>AE_OR2</type>
<position>390.5,-78</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>631 </input>
<output>
<ID>OUT</ID>653 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>675</ID>
<type>AE_DFF_LOW</type>
<position>395,-85</position>
<input>
<ID>IN_0</ID>653 </input>
<output>
<ID>OUT_0</ID>636 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>676</ID>
<type>AA_AND2</type>
<position>397.5,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>636 </input>
<output>
<ID>OUT</ID>634 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>677</ID>
<type>AA_AND2</type>
<position>401.5,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>788 </input>
<output>
<ID>OUT</ID>635 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>678</ID>
<type>AE_OR2</type>
<position>399.5,-78</position>
<input>
<ID>IN_0</ID>635 </input>
<input>
<ID>IN_1</ID>634 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>679</ID>
<type>AE_DFF_LOW</type>
<position>404.5,-85</position>
<input>
<ID>IN_0</ID>652 </input>
<output>
<ID>OUT_0</ID>639 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>680</ID>
<type>AA_AND2</type>
<position>407,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>637 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>681</ID>
<type>AA_AND2</type>
<position>411,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>789 </input>
<output>
<ID>OUT</ID>638 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>682</ID>
<type>AE_OR2</type>
<position>409,-78</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>637 </input>
<output>
<ID>OUT</ID>654 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>683</ID>
<type>AE_DFF_LOW</type>
<position>413.5,-85</position>
<input>
<ID>IN_0</ID>654 </input>
<output>
<ID>OUT_0</ID>642 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>684</ID>
<type>AA_AND2</type>
<position>416,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>642 </input>
<output>
<ID>OUT</ID>640 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>685</ID>
<type>AA_AND2</type>
<position>420,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>641 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>686</ID>
<type>AE_OR2</type>
<position>418,-78</position>
<input>
<ID>IN_0</ID>641 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>655 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>687</ID>
<type>AE_DFF_LOW</type>
<position>422.5,-85</position>
<input>
<ID>IN_0</ID>655 </input>
<output>
<ID>OUT_0</ID>645 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>688</ID>
<type>AA_AND2</type>
<position>425,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>645 </input>
<output>
<ID>OUT</ID>643 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_AND2</type>
<position>429,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>791 </input>
<output>
<ID>OUT</ID>644 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_OR2</type>
<position>427,-78</position>
<input>
<ID>IN_0</ID>644 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>656 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>691</ID>
<type>AE_DFF_LOW</type>
<position>431.5,-85</position>
<input>
<ID>IN_0</ID>656 </input>
<output>
<ID>OUT_0</ID>648 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>692</ID>
<type>AA_AND2</type>
<position>434,-72</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>648 </input>
<output>
<ID>OUT</ID>646 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>693</ID>
<type>AA_AND2</type>
<position>438,-72</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>776 </input>
<output>
<ID>OUT</ID>647 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>694</ID>
<type>AE_OR2</type>
<position>436,-78</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>646 </input>
<output>
<ID>OUT</ID>657 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>AE_DFF_LOW</type>
<position>440.5,-85</position>
<input>
<ID>IN_0</ID>657 </input>
<output>
<ID>OUT_0</ID>808 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>696</ID>
<type>BB_CLOCK</type>
<position>164.5,0.5</position>
<output>
<ID>CLK</ID>665 </output>
<gparam>angle 90</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>698</ID>
<type>AA_AND2</type>
<position>171.5,-2.5</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>700 </input>
<output>
<ID>OUT</ID>663 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>699</ID>
<type>AA_AND4</type>
<position>281.5,-82.5</position>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>714 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>700</ID>
<type>AE_DFF_LOW</type>
<position>375.5,-25.5</position>
<input>
<ID>IN_0</ID>777 </input>
<output>
<ID>OUT_0</ID>670 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>701</ID>
<type>AA_AND2</type>
<position>378,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>666 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>702</ID>
<type>AA_AND2</type>
<position>459.5,-100</position>
<input>
<ID>IN_0</ID>703 </input>
<input>
<ID>IN_1</ID>705 </input>
<output>
<ID>OUT</ID>702 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>703</ID>
<type>AA_AND2</type>
<position>382,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>778 </input>
<output>
<ID>OUT</ID>667 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>704</ID>
<type>AE_OR2</type>
<position>380,-18.5</position>
<input>
<ID>IN_0</ID>667 </input>
<input>
<ID>IN_1</ID>666 </input>
<output>
<ID>OUT</ID>691 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>705</ID>
<type>AA_AND2</type>
<position>474.5,-115.5</position>
<input>
<ID>IN_0</ID>709 </input>
<input>
<ID>IN_1</ID>709 </input>
<output>
<ID>OUT</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>706</ID>
<type>AE_DFF_LOW</type>
<position>384.5,-25.5</position>
<input>
<ID>IN_0</ID>691 </input>
<output>
<ID>OUT_0</ID>673 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>707</ID>
<type>AE_SMALL_INVERTER</type>
<position>444.5,-103</position>
<input>
<ID>IN_0</ID>712 </input>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>708</ID>
<type>AA_AND2</type>
<position>387,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>673 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>AA_AND2</type>
<position>391,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>779 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>710</ID>
<type>AE_OR2</type>
<position>389,-18.5</position>
<input>
<ID>IN_0</ID>672 </input>
<input>
<ID>IN_1</ID>671 </input>
<output>
<ID>OUT</ID>693 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>711</ID>
<type>AE_DFF_LOW</type>
<position>393.5,-25.5</position>
<input>
<ID>IN_0</ID>693 </input>
<output>
<ID>OUT_0</ID>676 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>712</ID>
<type>AA_AND2</type>
<position>396,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>676 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>713</ID>
<type>AA_AND2</type>
<position>400,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>780 </input>
<output>
<ID>OUT</ID>675 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>714</ID>
<type>AE_OR2</type>
<position>398,-18.5</position>
<input>
<ID>IN_0</ID>675 </input>
<input>
<ID>IN_1</ID>674 </input>
<output>
<ID>OUT</ID>692 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>715</ID>
<type>AE_DFF_LOW</type>
<position>403,-25.5</position>
<input>
<ID>IN_0</ID>692 </input>
<output>
<ID>OUT_0</ID>679 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>716</ID>
<type>AA_AND2</type>
<position>405.5,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>679 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>717</ID>
<type>AA_AND2</type>
<position>409.5,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>781 </input>
<output>
<ID>OUT</ID>678 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>718</ID>
<type>AE_OR2</type>
<position>407.5,-18.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>677 </input>
<output>
<ID>OUT</ID>694 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>719</ID>
<type>AE_DFF_LOW</type>
<position>412,-25.5</position>
<input>
<ID>IN_0</ID>694 </input>
<output>
<ID>OUT_0</ID>682 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_AND2</type>
<position>414.5,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>682 </input>
<output>
<ID>OUT</ID>680 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>721</ID>
<type>AA_AND2</type>
<position>418.5,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>807 </input>
<output>
<ID>OUT</ID>681 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>722</ID>
<type>AE_OR2</type>
<position>416.5,-18.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>680 </input>
<output>
<ID>OUT</ID>695 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>723</ID>
<type>AE_DFF_LOW</type>
<position>421,-25.5</position>
<input>
<ID>IN_0</ID>695 </input>
<output>
<ID>OUT_0</ID>685 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>724</ID>
<type>AA_AND2</type>
<position>423.5,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>685 </input>
<output>
<ID>OUT</ID>683 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>725</ID>
<type>AA_AND2</type>
<position>427.5,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>783 </input>
<output>
<ID>OUT</ID>684 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>726</ID>
<type>AE_OR2</type>
<position>425.5,-18.5</position>
<input>
<ID>IN_0</ID>684 </input>
<input>
<ID>IN_1</ID>683 </input>
<output>
<ID>OUT</ID>696 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_DFF_LOW</type>
<position>430,-25.5</position>
<input>
<ID>IN_0</ID>696 </input>
<output>
<ID>OUT_0</ID>688 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>728</ID>
<type>AA_AND2</type>
<position>432.5,-12.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>688 </input>
<output>
<ID>OUT</ID>686 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>729</ID>
<type>AA_AND2</type>
<position>436.5,-12.5</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>784 </input>
<output>
<ID>OUT</ID>687 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>730</ID>
<type>AE_OR2</type>
<position>434.5,-18.5</position>
<input>
<ID>IN_0</ID>687 </input>
<input>
<ID>IN_1</ID>686 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>731</ID>
<type>AE_DFF_LOW</type>
<position>439,-25.5</position>
<input>
<ID>IN_0</ID>697 </input>
<output>
<ID>OUT_0</ID>809 </output>
<input>
<ID>clock</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>732</ID>
<type>AE_SMALL_INVERTER</type>
<position>444.5,-107</position>
<input>
<ID>IN_0</ID>710 </input>
<output>
<ID>OUT_0</ID>690 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>733</ID>
<type>AE_OR2</type>
<position>467,-111.5</position>
<input>
<ID>IN_0</ID>709 </input>
<input>
<ID>IN_1</ID>698 </input>
<output>
<ID>OUT</ID>699 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>734</ID>
<type>AE_SMALL_INVERTER</type>
<position>459,-120</position>
<input>
<ID>IN_0</ID>690 </input>
<output>
<ID>OUT_0</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>735</ID>
<type>BB_CLOCK</type>
<position>449,-117.5</position>
<output>
<ID>CLK</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>736</ID>
<type>AA_AND2</type>
<position>461.5,-115.5</position>
<input>
<ID>IN_0</ID>689 </input>
<input>
<ID>IN_1</ID>668 </input>
<output>
<ID>OUT</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>737</ID>
<type>AA_REGISTER4</type>
<position>460,-107.5</position>
<output>
<ID>OUT_0</ID>705 </output>
<output>
<ID>OUT_3</ID>703 </output>
<input>
<ID>clear</ID>702 </input>
<input>
<ID>clock</ID>699 </input>
<input>
<ID>count_enable</ID>701 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>738</ID>
<type>AA_TOGGLE</type>
<position>453,-107.5</position>
<output>
<ID>OUT_0</ID>701 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>739</ID>
<type>AE_SMALL_INVERTER</type>
<position>450,-112.5</position>
<input>
<ID>IN_0</ID>702 </input>
<output>
<ID>OUT_0</ID>669 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>740</ID>
<type>AA_AND2</type>
<position>455,-113.5</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>690 </input>
<output>
<ID>OUT</ID>689 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>742</ID>
<type>AE_DFF_LOW</type>
<position>485.5,-102.5</position>
<input>
<ID>IN_0</ID>739 </input>
<output>
<ID>OUT_0</ID>720 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>743</ID>
<type>AA_AND2</type>
<position>488.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>720 </input>
<output>
<ID>OUT</ID>716 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>744</ID>
<type>AA_AND2</type>
<position>492.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>793 </input>
<output>
<ID>OUT</ID>717 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>745</ID>
<type>AE_OR2</type>
<position>490.5,-95.5</position>
<input>
<ID>IN_0</ID>717 </input>
<input>
<ID>IN_1</ID>716 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>746</ID>
<type>AA_AND4</type>
<position>281.5,-90.5</position>
<input>
<ID>IN_1</ID>798 </input>
<input>
<ID>IN_2</ID>719 </input>
<input>
<ID>IN_3</ID>796 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>AA_AND2</type>
<position>474,-92.5</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>711 </input>
<output>
<ID>OUT</ID>718 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>748</ID>
<type>AE_DFF_LOW</type>
<position>495.5,-102.5</position>
<input>
<ID>IN_0</ID>741 </input>
<output>
<ID>OUT_0</ID>723 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>749</ID>
<type>AA_AND2</type>
<position>498.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>723 </input>
<output>
<ID>OUT</ID>721 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>750</ID>
<type>AA_AND2</type>
<position>502.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>753 </input>
<output>
<ID>OUT</ID>722 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>751</ID>
<type>AE_OR2</type>
<position>500.5,-95.5</position>
<input>
<ID>IN_0</ID>722 </input>
<input>
<ID>IN_1</ID>721 </input>
<output>
<ID>OUT</ID>743 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>752</ID>
<type>AE_DFF_LOW</type>
<position>505.5,-102.5</position>
<input>
<ID>IN_0</ID>743 </input>
<output>
<ID>OUT_0</ID>726 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>753</ID>
<type>AA_AND2</type>
<position>508.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>726 </input>
<output>
<ID>OUT</ID>724 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>754</ID>
<type>AA_AND2</type>
<position>512.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>752 </input>
<output>
<ID>OUT</ID>725 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_OR2</type>
<position>510.5,-95.5</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>724 </input>
<output>
<ID>OUT</ID>742 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>756</ID>
<type>AE_DFF_LOW</type>
<position>515.5,-102.5</position>
<input>
<ID>IN_0</ID>742 </input>
<output>
<ID>OUT_0</ID>729 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>757</ID>
<type>AA_AND2</type>
<position>518.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>729 </input>
<output>
<ID>OUT</ID>727 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>AA_AND2</type>
<position>522.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>751 </input>
<output>
<ID>OUT</ID>728 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>759</ID>
<type>AE_OR2</type>
<position>520.5,-95.5</position>
<input>
<ID>IN_0</ID>728 </input>
<input>
<ID>IN_1</ID>727 </input>
<output>
<ID>OUT</ID>744 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>760</ID>
<type>AE_DFF_LOW</type>
<position>525.5,-102.5</position>
<input>
<ID>IN_0</ID>744 </input>
<output>
<ID>OUT_0</ID>732 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_AND2</type>
<position>528.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>732 </input>
<output>
<ID>OUT</ID>730 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>762</ID>
<type>AA_AND2</type>
<position>532.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>750 </input>
<output>
<ID>OUT</ID>731 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>763</ID>
<type>AE_OR2</type>
<position>530.5,-95.5</position>
<input>
<ID>IN_0</ID>731 </input>
<input>
<ID>IN_1</ID>730 </input>
<output>
<ID>OUT</ID>745 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>764</ID>
<type>AE_DFF_LOW</type>
<position>535.5,-102.5</position>
<input>
<ID>IN_0</ID>745 </input>
<output>
<ID>OUT_0</ID>735 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>765</ID>
<type>AA_AND2</type>
<position>538.5,-89.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>735 </input>
<output>
<ID>OUT</ID>733 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>766</ID>
<type>AA_AND2</type>
<position>542.5,-89.5</position>
<input>
<ID>IN_0</ID>775 </input>
<input>
<ID>IN_1</ID>749 </input>
<output>
<ID>OUT</ID>734 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>767</ID>
<type>AE_OR2</type>
<position>540.5,-95.5</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>733 </input>
<output>
<ID>OUT</ID>746 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>768</ID>
<type>AE_DFF_LOW</type>
<position>545.5,-102.5</position>
<input>
<ID>IN_0</ID>746 </input>
<output>
<ID>OUT_0</ID>738 </output>
<input>
<ID>clock</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>769</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579.5,-37.5,579.5,-30.5</points>
<intersection>-37.5 5</intersection>
<intersection>-30.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>579.5,-37.5,583.5,-37.5</points>
<connection>
<GID>785</GID>
<name>IN_4</name></connection>
<intersection>579.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>571.5,-30.5,579.5,-30.5</points>
<intersection>571.5 8</intersection>
<intersection>579.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>571.5,-31.5,571.5,-29.5</points>
<connection>
<GID>790</GID>
<name>OUT_0</name></connection>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<intersection>-30.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>770</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-23.5,571.5,-21.5</points>
<connection>
<GID>791</GID>
<name>OUT_0</name></connection>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>571.5,-22.5,580.5,-22.5</points>
<intersection>571.5 0</intersection>
<intersection>580.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>580.5,-36.5,580.5,-22.5</points>
<intersection>-36.5 5</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>580.5,-36.5,583.5,-36.5</points>
<connection>
<GID>785</GID>
<name>IN_5</name></connection>
<intersection>580.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,13,-22,39</points>
<connection>
<GID>55</GID>
<name>A_greater_B</name></connection>
<intersection>13 8</intersection>
<intersection>19 10</intersection>
<intersection>29 9</intersection>
<intersection>35 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-22,35,-17,35</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-22,13,-17,13</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-22,29,-21,29</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-22,19,-21,19</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>771</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-15.5,571.5,-13.5</points>
<connection>
<GID>792</GID>
<name>OUT_0</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>571.5,-14.5,581.5,-14.5</points>
<intersection>571.5 0</intersection>
<intersection>581.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>581.5,-35.5,581.5,-14.5</points>
<intersection>-35.5 5</intersection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>581.5,-35.5,583.5,-35.5</points>
<connection>
<GID>785</GID>
<name>IN_6</name></connection>
<intersection>581.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>772</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-7.5,571.5,-6.5</points>
<connection>
<GID>793</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571.5,-6.5,582.5,-6.5</points>
<intersection>571.5 0</intersection>
<intersection>582.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>582.5,-34.5,582.5,-6.5</points>
<intersection>-34.5 3</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>582.5,-34.5,583.5,-34.5</points>
<connection>
<GID>785</GID>
<name>IN_7</name></connection>
<intersection>582.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>773</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>586.5,-32.5,586.5,-32.5</points>
<connection>
<GID>785</GID>
<name>load</name></connection>
<connection>
<GID>794</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>774</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>559.5,-100.5,559.5,-72.5</points>
<intersection>-100.5 5</intersection>
<intersection>-72.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>558.5,-100.5,559.5,-100.5</points>
<connection>
<GID>772</GID>
<name>OUT_0</name></connection>
<intersection>559.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>559.5,-72.5,560.5,-72.5</points>
<connection>
<GID>661</GID>
<name>IN_0</name></connection>
<intersection>559.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>775</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-86.5,493.5,-85.5</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>482.5,-85.5,553.5,-85.5</points>
<connection>
<GID>799</GID>
<name>OUT_0</name></connection>
<intersection>493.5 0</intersection>
<intersection>503.5 5</intersection>
<intersection>513.5 6</intersection>
<intersection>523.5 7</intersection>
<intersection>533.5 8</intersection>
<intersection>543.5 10</intersection>
<intersection>553.5 11</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>503.5,-86.5,503.5,-85.5</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>513.5,-86.5,513.5,-85.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>523.5,-86.5,523.5,-85.5</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>533.5,-86.5,533.5,-85.5</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>543.5,-86.5,543.5,-85.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>553.5,-86.5,553.5,-85.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>-85.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-69,437,-58</points>
<connection>
<GID>693</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>355,-58,437,-58</points>
<intersection>355 2</intersection>
<intersection>437 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>355,-81.5,355,-58</points>
<intersection>-81.5 3</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>344,-81.5,355,-81.5</points>
<connection>
<GID>632</GID>
<name>OUT_7</name></connection>
<intersection>355 2</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361,-23.5,361,-5.5</points>
<intersection>-23.5 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-23.5,372.5,-23.5</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>361 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-5.5,361,-5.5</points>
<connection>
<GID>621</GID>
<name>OUT_0</name></connection>
<intersection>361 0</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381,-9.5,381,-4.5</points>
<connection>
<GID>703</GID>
<name>IN_1</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-4.5,381,-4.5</points>
<connection>
<GID>621</GID>
<name>OUT_1</name></connection>
<intersection>381 0</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>390,-9.5,390,-3.5</points>
<connection>
<GID>709</GID>
<name>IN_1</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-3.5,390,-3.5</points>
<connection>
<GID>621</GID>
<name>OUT_2</name></connection>
<intersection>390 0</intersection></hsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,-9.5,399,-2.5</points>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-2.5,399,-2.5</points>
<connection>
<GID>621</GID>
<name>OUT_3</name></connection>
<intersection>399 0</intersection></hsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>408.5,-9.5,408.5,-1.5</points>
<connection>
<GID>717</GID>
<name>IN_1</name></connection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-1.5,408.5,-1.5</points>
<connection>
<GID>621</GID>
<name>OUT_4</name></connection>
<intersection>408.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>370.5,-67.5,370.5,32.5</points>
<intersection>-67.5 59</intersection>
<intersection>-7.5 37</intersection>
<intersection>32.5 35</intersection></vsegment>
<vsegment>
<ID>22</ID>
<points>252,-30.5,252,32.5</points>
<intersection>-30.5 88</intersection>
<intersection>32.5 35</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>252,32.5,370.5,32.5</points>
<intersection>252 22</intersection>
<intersection>370.5 2</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>370.5,-7.5,433.5,-7.5</points>
<intersection>370.5 2</intersection>
<intersection>379 80</intersection>
<intersection>388 52</intersection>
<intersection>397 53</intersection>
<intersection>406.5 54</intersection>
<intersection>415.5 55</intersection>
<intersection>424.5 56</intersection>
<intersection>433.5 51</intersection></hsegment>
<vsegment>
<ID>51</ID>
<points>433.5,-9.5,433.5,-7.5</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<vsegment>
<ID>52</ID>
<points>388,-9.5,388,-7.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<vsegment>
<ID>53</ID>
<points>397,-9.5,397,-7.5</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>406.5,-9.5,406.5,-7.5</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<vsegment>
<ID>55</ID>
<points>415.5,-9.5,415.5,-7.5</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<vsegment>
<ID>56</ID>
<points>424.5,-9.5,424.5,-7.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<hsegment>
<ID>59</ID>
<points>370.5,-67.5,435,-67.5</points>
<intersection>370.5 2</intersection>
<intersection>380.5 60</intersection>
<intersection>389.5 74</intersection>
<intersection>398.5 75</intersection>
<intersection>408 76</intersection>
<intersection>417 77</intersection>
<intersection>426 78</intersection>
<intersection>435 73</intersection></hsegment>
<vsegment>
<ID>60</ID>
<points>380.5,-69,380.5,-67.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>435,-69,435,-67.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>389.5,-69,389.5,-67.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>398.5,-69,398.5,-67.5</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>408,-69,408,-67.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>417,-69,417,-67.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>426,-69,426,-67.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-67.5 59</intersection></vsegment>
<vsegment>
<ID>80</ID>
<points>379,-9.5,379,-7.5</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>-7.5 37</intersection></vsegment>
<hsegment>
<ID>88</ID>
<points>208,-30.5,252,-30.5</points>
<connection>
<GID>669</GID>
<name>OUT</name></connection>
<intersection>252 22</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-9.5,426.5,0.5</points>
<connection>
<GID>725</GID>
<name>IN_1</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,0.5,426.5,0.5</points>
<connection>
<GID>621</GID>
<name>OUT_6</name></connection>
<intersection>426.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>435.5,-9.5,435.5,1.5</points>
<connection>
<GID>729</GID>
<name>IN_1</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,1.5,435.5,1.5</points>
<connection>
<GID>621</GID>
<name>OUT_7</name></connection>
<intersection>435.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>785</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-88.5,362,-83</points>
<intersection>-88.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344,-88.5,362,-88.5</points>
<connection>
<GID>632</GID>
<name>OUT_0</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>362,-83,374,-83</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>382.5,-69,382.5,-64</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361,-64,382.5,-64</points>
<intersection>361 2</intersection>
<intersection>382.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>361,-87.5,361,-64</points>
<intersection>-87.5 5</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>344,-87.5,361,-87.5</points>
<connection>
<GID>632</GID>
<name>OUT_1</name></connection>
<intersection>361 2</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>391.5,-69,391.5,-63</points>
<connection>
<GID>673</GID>
<name>IN_1</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>360,-63,391.5,-63</points>
<intersection>360 2</intersection>
<intersection>391.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>360,-86.5,360,-63</points>
<intersection>-86.5 3</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>344,-86.5,360,-86.5</points>
<connection>
<GID>632</GID>
<name>OUT_2</name></connection>
<intersection>360 2</intersection></hsegment></shape></wire>
<wire>
<ID>788</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-69,400.5,-62</points>
<connection>
<GID>677</GID>
<name>IN_1</name></connection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-62,400.5,-62</points>
<intersection>359 2</intersection>
<intersection>400.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>359,-85.5,359,-62</points>
<intersection>-85.5 3</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>344,-85.5,359,-85.5</points>
<connection>
<GID>632</GID>
<name>OUT_3</name></connection>
<intersection>359 2</intersection></hsegment></shape></wire>
<wire>
<ID>789</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410,-69,410,-61</points>
<connection>
<GID>681</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>358,-61,410,-61</points>
<intersection>358 2</intersection>
<intersection>410 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>358,-84.5,358,-61</points>
<intersection>-84.5 3</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>344,-84.5,358,-84.5</points>
<connection>
<GID>632</GID>
<name>OUT_4</name></connection>
<intersection>358 2</intersection></hsegment></shape></wire>
<wire>
<ID>790</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,-69,419,-60</points>
<connection>
<GID>685</GID>
<name>IN_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-60,419,-60</points>
<intersection>357 2</intersection>
<intersection>419 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>357,-83.5,357,-60</points>
<intersection>-83.5 5</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>344,-83.5,357,-83.5</points>
<connection>
<GID>632</GID>
<name>OUT_5</name></connection>
<intersection>357 2</intersection></hsegment></shape></wire>
<wire>
<ID>791</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>428,-69,428,-59</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356,-59,428,-59</points>
<intersection>356 2</intersection>
<intersection>428 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>356,-82.5,356,-59</points>
<intersection>-82.5 3</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>344,-82.5,356,-82.5</points>
<connection>
<GID>632</GID>
<name>OUT_6</name></connection>
<intersection>356 2</intersection></hsegment></shape></wire>
<wire>
<ID>792</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>578.5,-108,578.5,-13.5</points>
<intersection>-108 1</intersection>
<intersection>-69.5 4</intersection>
<intersection>-61.5 3</intersection>
<intersection>-53.5 10</intersection>
<intersection>-48.5 31</intersection>
<intersection>-45.5 9</intersection>
<intersection>-37.5 8</intersection>
<intersection>-29.5 11</intersection>
<intersection>-21.5 12</intersection>
<intersection>-13.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>570.5,-108,578.5,-108</points>
<connection>
<GID>810</GID>
<name>OUT</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>574.5,-61.5,578.5,-61.5</points>
<connection>
<GID>787</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>574.5,-69.5,578.5,-69.5</points>
<connection>
<GID>786</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>574.5,-13.5,578.5,-13.5</points>
<connection>
<GID>793</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>574.5,-37.5,578.5,-37.5</points>
<connection>
<GID>790</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>574.5,-45.5,578.5,-45.5</points>
<connection>
<GID>789</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>574.5,-53.5,578.5,-53.5</points>
<connection>
<GID>788</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>574.5,-29.5,578.5,-29.5</points>
<connection>
<GID>791</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>574.5,-21.5,578.5,-21.5</points>
<connection>
<GID>792</GID>
<name>clock</name></connection>
<intersection>578.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>578.5,-48.5,586.5,-48.5</points>
<intersection>578.5 0</intersection>
<intersection>586.5 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>586.5,-48.5,586.5,-47.5</points>
<connection>
<GID>795</GID>
<name>IN_0</name></connection>
<intersection>-48.5 31</intersection></vsegment></shape></wire>
<wire>
<ID>793</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>491.5,-86.5,491.5,-82</points>
<connection>
<GID>744</GID>
<name>IN_1</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-82,491.5,-82</points>
<connection>
<GID>774</GID>
<name>OUT_1</name></connection>
<intersection>491.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>794</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>586.5,-43.5,586.5,-43.5</points>
<connection>
<GID>785</GID>
<name>clock</name></connection>
<connection>
<GID>795</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,7,73,15.5</points>
<intersection>7 2</intersection>
<intersection>15.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67,7,73,7</points>
<intersection>67 3</intersection>
<intersection>73 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,7,67,8</points>
<connection>
<GID>39</GID>
<name>A_greater_B</name></connection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>73,15.5,75,15.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>795</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>141,-20,141,-4.5</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>-13 10</intersection>
<intersection>-4.5 31</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>141,-13,144.5,-13</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<intersection>141 7</intersection>
<intersection>144 32</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>141,-4.5,146,-4.5</points>
<connection>
<GID>655</GID>
<name>OUT</name></connection>
<intersection>141 7</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>144,-13,144,-11</points>
<intersection>-13 10</intersection>
<intersection>-11 33</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>144,-11,148.5,-11</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>144 32</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-11,74,14.5</points>
<intersection>-11 2</intersection>
<intersection>14.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67,-11,74,-11</points>
<intersection>67 3</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-11,67,-10</points>
<connection>
<GID>49</GID>
<name>A_greater_B</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>74,14.5,75,14.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>796</ID>
<shape>
<vsegment>
<ID>21</ID>
<points>276.5,-109.5,276.5,42</points>
<intersection>-109.5 33</intersection>
<intersection>-93.5 27</intersection>
<intersection>-77.5 26</intersection>
<intersection>-61.5 25</intersection>
<intersection>-35 68</intersection>
<intersection>-19 62</intersection>
<intersection>-3 61</intersection>
<intersection>13 60</intersection>
<intersection>42 55</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>276.5,-61.5,278.5,-61.5</points>
<connection>
<GID>612</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>276.5,-77.5,278.5,-77.5</points>
<connection>
<GID>658</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>276.5,-93.5,278.5,-93.5</points>
<connection>
<GID>746</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>276.5,-109.5,278.5,-109.5</points>
<connection>
<GID>806</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>55</ID>
<points>143.5,42,454.5,42</points>
<connection>
<GID>805</GID>
<name>OUT_0</name></connection>
<intersection>276.5 21</intersection>
<intersection>277.5 70</intersection>
<intersection>454.5 66</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>276.5,13,278.5,13</points>
<connection>
<GID>558</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>61</ID>
<points>276.5,-3,278.5,-3</points>
<connection>
<GID>562</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>276.5,-19,278.5,-19</points>
<connection>
<GID>566</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<vsegment>
<ID>66</ID>
<points>454.5,-52,454.5,42</points>
<connection>
<GID>660</GID>
<name>SEL_0</name></connection>
<intersection>42 55</intersection></vsegment>
<hsegment>
<ID>68</ID>
<points>276.5,-35,278.5,-35</points>
<connection>
<GID>570</GID>
<name>IN_3</name></connection>
<intersection>276.5 21</intersection></hsegment>
<vsegment>
<ID>70</ID>
<points>277.5,37,277.5,42</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<intersection>42 55</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,16.5,74,25</points>
<intersection>16.5 6</intersection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67,25,74,25</points>
<intersection>67 3</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,25,67,26</points>
<connection>
<GID>54</GID>
<name>A_greater_B</name></connection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>74,16.5,75,16.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>797</ID>
<shape>
<vsegment>
<ID>24</ID>
<points>274.5,-107.5,274.5,40</points>
<intersection>-107.5 39</intersection>
<intersection>-99.5 32</intersection>
<intersection>-75.5 30</intersection>
<intersection>-67.5 28</intersection>
<intersection>-33 80</intersection>
<intersection>-25 73</intersection>
<intersection>-1 71</intersection>
<intersection>7 69</intersection>
<intersection>40 64</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>274.5,-67.5,278.5,-67.5</points>
<connection>
<GID>630</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>274.5,-75.5,278.5,-75.5</points>
<connection>
<GID>658</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>274.5,-99.5,278.5,-99.5</points>
<connection>
<GID>800</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>274.5,-107.5,278.5,-107.5</points>
<connection>
<GID>806</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>64</ID>
<points>143.5,40,453.5,40</points>
<connection>
<GID>804</GID>
<name>OUT_0</name></connection>
<intersection>274.5 24</intersection>
<intersection>275.5 77</intersection>
<intersection>453.5 78</intersection></hsegment>
<hsegment>
<ID>69</ID>
<points>274.5,7,278.5,7</points>
<connection>
<GID>560</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>274.5,-1,278.5,-1</points>
<connection>
<GID>562</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<hsegment>
<ID>73</ID>
<points>274.5,-25,278.5,-25</points>
<connection>
<GID>568</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment>
<vsegment>
<ID>77</ID>
<points>275.5,37,275.5,40</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>40 64</intersection></vsegment>
<vsegment>
<ID>78</ID>
<points>453.5,-52,453.5,40</points>
<connection>
<GID>660</GID>
<name>SEL_1</name></connection>
<intersection>40 64</intersection></vsegment>
<hsegment>
<ID>80</ID>
<points>274.5,-33,278.5,-33</points>
<connection>
<GID>570</GID>
<name>IN_2</name></connection>
<intersection>274.5 24</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,20.5,78,22.5</points>
<connection>
<GID>56</GID>
<name>load</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>798</ID>
<shape>
<vsegment>
<ID>23</ID>
<points>272.5,-105.5,272.5,38</points>
<intersection>-105.5 39</intersection>
<intersection>-97.5 31</intersection>
<intersection>-89.5 29</intersection>
<intersection>-81.5 27</intersection>
<intersection>-31 80</intersection>
<intersection>-23 72</intersection>
<intersection>-15 70</intersection>
<intersection>-7 68</intersection>
<intersection>38 63</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>272.5,-81.5,278.5,-81.5</points>
<connection>
<GID>699</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>272.5,-89.5,278.5,-89.5</points>
<connection>
<GID>746</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>272.5,-97.5,278.5,-97.5</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>272.5,-105.5,278.5,-105.5</points>
<connection>
<GID>806</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>63</ID>
<points>143.5,38,452.5,38</points>
<connection>
<GID>803</GID>
<name>OUT_0</name></connection>
<intersection>272.5 23</intersection>
<intersection>273.5 87</intersection>
<intersection>452.5 78</intersection></hsegment>
<hsegment>
<ID>68</ID>
<points>272.5,-7,278.5,-7</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>70</ID>
<points>272.5,-15,278.5,-15</points>
<connection>
<GID>566</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<hsegment>
<ID>72</ID>
<points>272.5,-23,278.5,-23</points>
<connection>
<GID>568</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<vsegment>
<ID>78</ID>
<points>452.5,-52,452.5,38</points>
<connection>
<GID>660</GID>
<name>SEL_2</name></connection>
<intersection>38 63</intersection></vsegment>
<hsegment>
<ID>80</ID>
<points>272.5,-31,278.5,-31</points>
<connection>
<GID>570</GID>
<name>IN_1</name></connection>
<intersection>272.5 23</intersection></hsegment>
<vsegment>
<ID>87</ID>
<points>273.5,37,273.5,38</points>
<connection>
<GID>572</GID>
<name>IN_0</name></connection>
<intersection>38 63</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,9.5,78,11.5</points>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>799</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319,-50.5,319,23.5</points>
<intersection>-50.5 26</intersection>
<intersection>-39 1</intersection>
<intersection>-31.5 8</intersection>
<intersection>-23 7</intersection>
<intersection>-14.5 9</intersection>
<intersection>-6.5 14</intersection>
<intersection>1 13</intersection>
<intersection>8.5 12</intersection>
<intersection>16 11</intersection>
<intersection>23.5 10</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319,-39,337,-39</points>
<intersection>319 0</intersection>
<intersection>337 16</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>312,-23,319,-23</points>
<connection>
<GID>623</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>312,-31.5,319,-31.5</points>
<connection>
<GID>622</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>312,-14.5,319,-14.5</points>
<connection>
<GID>624</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>312,23.5,319,23.5</points>
<connection>
<GID>629</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>312,16,319,16</points>
<connection>
<GID>628</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>312,8.5,319,8.5</points>
<connection>
<GID>627</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>312,1,319,1</points>
<connection>
<GID>626</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>312,-6.5,319,-6.5</points>
<connection>
<GID>625</GID>
<name>clock</name></connection>
<intersection>319 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>337,-39,337,-11.5</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>284.5,-50.5,319,-50.5</points>
<connection>
<GID>575</GID>
<name>OUT</name></connection>
<intersection>319 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-34,32,-33,32</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<connection>
<GID>77</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>800</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>322.5,-115.5,322.5,-58</points>
<intersection>-115.5 4</intersection>
<intersection>-106 11</intersection>
<intersection>-98 12</intersection>
<intersection>-90 9</intersection>
<intersection>-82 8</intersection>
<intersection>-74 7</intersection>
<intersection>-66 6</intersection>
<intersection>-58 50</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>285.5,-115.5,339,-115.5</points>
<intersection>285.5 48</intersection>
<intersection>314 52</intersection>
<intersection>322.5 0</intersection>
<intersection>339 39</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>314,-66,322.5,-66</points>
<connection>
<GID>639</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>314,-74,322.5,-74</points>
<connection>
<GID>638</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>314,-82,322.5,-82</points>
<connection>
<GID>637</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>314,-90,322.5,-90</points>
<connection>
<GID>636</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>314,-106,322.5,-106</points>
<connection>
<GID>634</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>314,-98,322.5,-98</points>
<connection>
<GID>635</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<vsegment>
<ID>39</ID>
<points>339,-115.5,339,-94.5</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-115.5 4</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>285.5,-115.5,285.5,-58.5</points>
<intersection>-115.5 4</intersection>
<intersection>-58.5 51</intersection></vsegment>
<hsegment>
<ID>50</ID>
<points>314,-58,322.5,-58</points>
<connection>
<GID>640</GID>
<name>clock</name></connection>
<intersection>322.5 0</intersection></hsegment>
<hsegment>
<ID>51</ID>
<points>284.5,-58.5,285.5,-58.5</points>
<connection>
<GID>612</GID>
<name>OUT</name></connection>
<intersection>285.5 48</intersection></hsegment>
<vsegment>
<ID>52</ID>
<points>314,-115.5,314,-114.5</points>
<connection>
<GID>633</GID>
<name>clock</name></connection>
<intersection>-115.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-31,32,-30,32</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>801</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,33.5,147.5,33.5</points>
<connection>
<GID>811</GID>
<name>IN_0</name></connection>
<connection>
<GID>853</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-41,32,-40,32</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>75</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>802</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>145.5,22,145.5,30.5</points>
<connection>
<GID>812</GID>
<name>CLK</name></connection>
<intersection>22 5</intersection>
<intersection>30.5 7</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>145.5,22,147.5,22</points>
<connection>
<GID>813</GID>
<name>clock</name></connection>
<intersection>145.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>145.5,30.5,147.5,30.5</points>
<connection>
<GID>811</GID>
<name>clock</name></connection>
<intersection>145.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-44,32,-43,32</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>73</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>803</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,25,147.5,25</points>
<connection>
<GID>813</GID>
<name>IN_0</name></connection>
<connection>
<GID>854</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-51,32,-50,32</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>804</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-13,148.5,-13</points>
<connection>
<GID>814</GID>
<name>OUT_0</name></connection>
<connection>
<GID>815</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-54,32,-53,32</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>805</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>337,-7.5,337,-7.5</points>
<connection>
<GID>552</GID>
<name>OUT_0</name></connection>
<connection>
<GID>621</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-61,32,-60,32</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>806</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>339,-90.5,339,-90.5</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<connection>
<GID>632</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>807</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>417.5,-9.5,417.5,-0.5</points>
<connection>
<GID>721</GID>
<name>IN_1</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-0.5,417.5,-0.5</points>
<connection>
<GID>621</GID>
<name>OUT_5</name></connection>
<intersection>417.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-64,32,-63,32</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>808</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,-83,444.5,-60</points>
<intersection>-83 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>443.5,-83,444.5,-83</points>
<connection>
<GID>695</GID>
<name>OUT_0</name></connection>
<intersection>444.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444.5,-60,450.5,-60</points>
<connection>
<GID>660</GID>
<name>IN_1</name></connection>
<intersection>444.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,24,-62,26</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,24,-60,24</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>809</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,-61,444,-23.5</points>
<intersection>-61 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>442,-23.5,444,-23.5</points>
<connection>
<GID>731</GID>
<name>OUT_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,-61,450.5,-61</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-31,38,-31,38</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-41,38,-41,38</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>810</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>155,44,562.5,44</points>
<intersection>155 13</intersection>
<intersection>458.5 24</intersection>
<intersection>562.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>562.5,-69,562.5,44</points>
<connection>
<GID>661</GID>
<name>SEL_0</name></connection>
<intersection>44 7</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>155,-5.5,155,44</points>
<intersection>-5.5 14</intersection>
<intersection>33.5 35</intersection>
<intersection>44 7</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>152,-5.5,173.5,-5.5</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<intersection>155 13</intersection>
<intersection>173.5 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>173.5,-45.5,173.5,-5.5</points>
<intersection>-45.5 19</intersection>
<intersection>-29.5 22</intersection>
<intersection>-5.5 14</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>173.5,-45.5,175,-45.5</points>
<connection>
<GID>656</GID>
<name>IN_1</name></connection>
<intersection>173.5 18</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>173.5,-29.5,184.5,-29.5</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>173.5 18</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>458.5,-82.5,458.5,44</points>
<intersection>-82.5 31</intersection>
<intersection>44 7</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>457,-82.5,458.5,-82.5</points>
<connection>
<GID>809</GID>
<name>IN_0</name></connection>
<intersection>458.5 24</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>153.5,33.5,155,33.5</points>
<connection>
<GID>811</GID>
<name>OUT_0</name></connection>
<intersection>155 13</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-51,38,-51,38</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>811</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287.5,-31.5,287.5,24</points>
<intersection>-31.5 2</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,24,287.5,24</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<intersection>287.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>287.5,-31.5,309,-31.5</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>287.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-61,38,-61,38</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>812</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-114.5,286.5,16</points>
<intersection>-114.5 2</intersection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,16,286.5,16</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>286.5,-114.5,311,-114.5</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,26.5,-57,38</points>
<intersection>26.5 1</intersection>
<intersection>38 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,26.5,-54,26.5</points>
<intersection>-57 0</intersection>
<intersection>-54 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-54,24,-54,26.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-57,38,-55,38</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,26.5,-47,38</points>
<intersection>26.5 1</intersection>
<intersection>38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,26.5,-44,26.5</points>
<intersection>-47 0</intersection>
<intersection>-44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,38,-45,38</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44,24,-44,26.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,26.5,-37,38</points>
<intersection>26.5 1</intersection>
<intersection>38 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,26.5,-34,26.5</points>
<intersection>-37 0</intersection>
<intersection>-34 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34,24,-34,26.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-37,38,-35,38</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,38,-63,44</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,44,-31,44</points>
<intersection>-68 16</intersection>
<intersection>-63 0</intersection>
<intersection>-61 3</intersection>
<intersection>-53 5</intersection>
<intersection>-51 7</intersection>
<intersection>-43 9</intersection>
<intersection>-41 11</intersection>
<intersection>-33 13</intersection>
<intersection>-31 15</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-61,42,-61,44</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-53,38,-53,44</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-51,42,-51,44</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-43,38,-43,44</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-41,42,-41,44</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-33,38,-33,44</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>-31,42,-31,44</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>44 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>-68,9,-68,44</points>
<intersection>9 17</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-73,9,-31,9</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-68 16</intersection>
<intersection>-63 39</intersection>
<intersection>-61 22</intersection>
<intersection>-53 35</intersection>
<intersection>-51 26</intersection>
<intersection>-43 36</intersection>
<intersection>-41 30</intersection>
<intersection>-33 37</intersection>
<intersection>-31 34</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-61,8,-61,9</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-51,8,-51,9</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-41,8,-41,9</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>-31,8,-31,9</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>35</ID>
<points>-53,4,-53,9</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>-43,4,-43,9</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>-33,4,-33,9</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>-63,4,-63,9</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>9 17</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,24,-52,26</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,24,-50,24</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,24,-42,26</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42,24,-40,24</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-42 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,24,-32,26</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,24,-30,24</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,85,-86,85</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<connection>
<GID>834</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-34,-2,-33,-2</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89,83,-89,84</points>
<intersection>83 2</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-89,84,-86,84</points>
<connection>
<GID>834</GID>
<name>IN_2</name></connection>
<intersection>-89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90,83,-89,83</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<intersection>-89 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-31,-2,-30,-2</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-41,-2,-40,-2</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,79,-87,82</points>
<intersection>79 2</intersection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,82,-86,82</points>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90,79,-87,79</points>
<connection>
<GID>409</GID>
<name>OUT_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-44,-2,-43,-2</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>95</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-51,-2,-50,-2</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>92</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-54,-2,-53,-2</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-61,-2,-60,-2</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-64,-2,-63,-2</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-10,-62,-8</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-10,-60,-10</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-31,4,-31,4</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-41,4,-41,4</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-51,4,-51,4</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-61,4,-61,4</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-7.5,-57,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,-7.5,-54,-7.5</points>
<intersection>-57 0</intersection>
<intersection>-54 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-54,-10,-54,-7.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-57,4,-55,4</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,-7.5,-47,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,-7.5,-44,-7.5</points>
<intersection>-47 0</intersection>
<intersection>-44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,4,-45,4</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44,-10,-44,-7.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-7.5,-37,4</points>
<intersection>-7.5 1</intersection>
<intersection>4 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,-7.5,-34,-7.5</points>
<intersection>-37 0</intersection>
<intersection>-34 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34,-10,-34,-7.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-37,4,-35,4</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,52,-86,52</points>
<connection>
<GID>836</GID>
<name>IN_7</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-10,-52,-8</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-10,-50,-10</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-52 0</intersection></hsegment></shape></wire>
<wire>
<ID>836</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93,50,-93,51</points>
<intersection>50 2</intersection>
<intersection>51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93,51,-86,51</points>
<connection>
<GID>836</GID>
<name>IN_6</name></connection>
<intersection>-93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-94,50,-93,50</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-93 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-10,-42,-8</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-42,-10,-40,-10</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-42 0</intersection></hsegment></shape></wire>
<wire>
<ID>837</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87,36,-87,45</points>
<intersection>36 2</intersection>
<intersection>45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87,45,-86,45</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<intersection>-87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-94,36,-87,36</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-87 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-10,-32,-8</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32,-10,-30,-10</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>838</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,38,-88,46</points>
<intersection>38 2</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-88,46,-86,46</points>
<connection>
<GID>836</GID>
<name>IN_1</name></connection>
<intersection>-88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-94,38,-88,38</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-88 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,4,-65,4</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>839</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89,40,-89,47</points>
<intersection>40 2</intersection>
<intersection>47 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-94,40,-89,40</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-89 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-89,47,-86,47</points>
<connection>
<GID>836</GID>
<name>IN_2</name></connection>
<intersection>-89 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-65,38,-65,38</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>840</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90,42,-90,48</points>
<intersection>42 2</intersection>
<intersection>48 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-94,42,-90,42</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-90 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-90,48,-86,48</points>
<connection>
<GID>836</GID>
<name>IN_3</name></connection>
<intersection>-90 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,29,-17,29</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>841</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91,46,-91,49</points>
<intersection>46 3</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91,49,-86,49</points>
<connection>
<GID>836</GID>
<name>IN_4</name></connection>
<intersection>-91 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-94,46,-91,46</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-91 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,23,47,23</points>
<connection>
<GID>53</GID>
<name>IN_B_3</name></connection>
<intersection>7 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7,23,7,33</points>
<intersection>23 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6,33,8,33</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>7 3</intersection></hsegment></shape></wire>
<wire>
<ID>842</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92,48,-92,50</points>
<intersection>48 2</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-92,50,-86,50</points>
<connection>
<GID>836</GID>
<name>IN_5</name></connection>
<intersection>-92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-94,48,-92,48</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-92 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,24,47,24</points>
<connection>
<GID>53</GID>
<name>IN_B_2</name></connection>
<intersection>15 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,24,15,33</points>
<intersection>24 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14,33,16,33</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>15 3</intersection></hsegment></shape></wire>
<wire>
<ID>843</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,52,-24,52</points>
<connection>
<GID>836</GID>
<name>OUT_7</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>-69 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-69,13,-69,52</points>
<intersection>13 4</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-69,13,-29,13</points>
<intersection>-69 3</intersection>
<intersection>-29 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-29,4,-29,13</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>13 4</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,25,47,25</points>
<connection>
<GID>53</GID>
<name>IN_B_1</name></connection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,25,23,33</points>
<intersection>25 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>22,33,24,33</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>23 3</intersection></hsegment></shape></wire>
<wire>
<ID>844</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,51,-24,51</points>
<connection>
<GID>836</GID>
<name>OUT_6</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>-70 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-70,12,-70,51</points>
<intersection>12 4</intersection>
<intersection>51 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-70,12,-39,12</points>
<intersection>-70 3</intersection>
<intersection>-39 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-39,4,-39,12</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>12 4</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2,33,0,33</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>845</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,50,-24,50</points>
<connection>
<GID>836</GID>
<name>OUT_5</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>-71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71,11,-71,50</points>
<intersection>11 4</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-71,11,-49,11</points>
<intersection>-71 3</intersection>
<intersection>-49 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-49,4,-49,11</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>11 4</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,17,8.5,17</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>7.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>7.5,9,7.5,17</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>17 1</intersection></vsegment></shape></wire>
<wire>
<ID>846</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,49,-24,49</points>
<connection>
<GID>836</GID>
<name>OUT_4</name></connection>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>-72 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-72,10,-72,49</points>
<intersection>10 4</intersection>
<intersection>49 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-72,10,-59,10</points>
<intersection>-72 3</intersection>
<intersection>-59 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-59,4,-59,10</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>10 4</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,17,16.5,17</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>15.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>15.5,9,15.5,17</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>17 1</intersection></vsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,38,-29,48</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82,48,-25,48</points>
<connection>
<GID>836</GID>
<name>OUT_3</name></connection>
<intersection>-29 0</intersection>
<intersection>-25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-25,45,-25,48</points>
<intersection>45 4</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-25,45,-24,45</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-25 3</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,17,24.5,17</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>23.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>23.5,9,23.5,17</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>17 1</intersection></vsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,44,-26,47</points>
<intersection>44 1</intersection>
<intersection>47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,44,-24,44</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,47,-26,47</points>
<connection>
<GID>836</GID>
<name>OUT_2</name></connection>
<intersection>-39 3</intersection>
<intersection>-26 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-39,38,-39,47</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>47 2</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-2,17,0,17</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<connection>
<GID>120</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,43,-27,46</points>
<intersection>43 1</intersection>
<intersection>46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,43,-24,43</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,46,-27,46</points>
<connection>
<GID>836</GID>
<name>OUT_1</name></connection>
<intersection>-49 3</intersection>
<intersection>-27 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-49,38,-49,46</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>46 2</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,24,-23,37</points>
<intersection>24 2</intersection>
<intersection>31 3</intersection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23,37,-17,37</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24,24,-23,24</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23,31,-17,31</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>850</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,42,-28,45</points>
<intersection>42 1</intersection>
<intersection>45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,42,-24,42</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-82,45,-28,45</points>
<connection>
<GID>836</GID>
<name>OUT_0</name></connection>
<intersection>-59 3</intersection>
<intersection>-28 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-59,38,-59,45</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>45 2</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,-10,-23,21</points>
<intersection>-10 2</intersection>
<intersection>15 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23,21,-17,21</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24,-10,-23,-10</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-23,15,-17,15</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,113,-88.5,113</points>
<intersection>-104.5 5</intersection>
<intersection>-88.5 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-104.5,81,-104.5,113</points>
<intersection>81 6</intersection>
<intersection>113 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-104.5,81,-93,81</points>
<connection>
<GID>848</GID>
<name>N_in0</name></connection>
<intersection>-104.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-88.5,113,-88.5,115</points>
<intersection>113 1</intersection>
<intersection>115 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-89.5,115,-87.5,115</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>-88.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,34,-10,36</points>
<intersection>34 1</intersection>
<intersection>36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,34,-8,34</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,36,-10,36</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>852</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88,81,-88,83</points>
<intersection>81 1</intersection>
<intersection>83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91,81,-88,81</points>
<connection>
<GID>848</GID>
<name>N_in1</name></connection>
<intersection>-88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88,83,-86,83</points>
<connection>
<GID>834</GID>
<name>IN_1</name></connection>
<intersection>-88 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,20,-10,32</points>
<intersection>20 2</intersection>
<intersection>32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,32,-8,32</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,20,-10,20</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>853</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-105.5,54.5,-105.5,118</points>
<intersection>54.5 7</intersection>
<intersection>87.5 3</intersection>
<intersection>118 11</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-122,87.5,-84,87.5</points>
<connection>
<GID>832</GID>
<name>OUT_0</name></connection>
<intersection>-105.5 0</intersection>
<intersection>-84 9</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-105.5,54.5,-84,54.5</points>
<intersection>-105.5 0</intersection>
<intersection>-84 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-84,53.5,-84,54.5</points>
<connection>
<GID>836</GID>
<name>ENABLE_0</name></connection>
<intersection>54.5 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-84,86.5,-84,87.5</points>
<connection>
<GID>834</GID>
<name>ENABLE_0</name></connection>
<intersection>87.5 3</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-105.5,118,-84.5,118</points>
<intersection>-105.5 0</intersection>
<intersection>-84.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-84.5,117,-84.5,118</points>
<connection>
<GID>846</GID>
<name>ENABLE_0</name></connection>
<intersection>118 11</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,18,-9,30</points>
<intersection>18 5</intersection>
<intersection>30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11,30,-9,30</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>-9 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-9,18,-8,18</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,33.5,126,33.5</points>
<connection>
<GID>801</GID>
<name>OUT_0</name></connection>
<connection>
<GID>853</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,14,-10,16</points>
<intersection>14 2</intersection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,16,-8,16</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,14,-10,14</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>855</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,25,126,25</points>
<connection>
<GID>854</GID>
<name>IN_0</name></connection>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,19,-17,19</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,9,31.5,17</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>17 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>30.5,17,31.5,17</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,107.5,175.5,111</points>
<connection>
<GID>444</GID>
<name>clock</name></connection>
<intersection>107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,107.5,175.5,107.5</points>
<connection>
<GID>446</GID>
<name>CLK</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,1,31.5,5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,125,126,125</points>
<connection>
<GID>443</GID>
<name>OUT_0</name></connection>
<connection>
<GID>857</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,1,30.5,4</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>4 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>23.5,4,23.5,5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,4,30.5,4</points>
<intersection>23.5 1</intersection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,131,126,131</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<connection>
<GID>856</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,1,29.5,3</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>3 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>15.5,3,15.5,5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15.5,3,29.5,3</points>
<intersection>15.5 1</intersection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,28,106,134</points>
<intersection>28 11</intersection>
<intersection>36.5 9</intersection>
<intersection>108.5 1</intersection>
<intersection>128 5</intersection>
<intersection>134 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,108.5,106,108.5</points>
<connection>
<GID>134</GID>
<name>N_in1</name></connection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>106,128,129,128</points>
<intersection>106 0</intersection>
<intersection>129 8</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>106,134,129,134</points>
<intersection>106 0</intersection>
<intersection>129 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>129,133,129,134</points>
<connection>
<GID>856</GID>
<name>ENABLE_0</name></connection>
<intersection>134 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>129,127,129,128</points>
<connection>
<GID>857</GID>
<name>ENABLE_0</name></connection>
<intersection>128 5</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>106,36.5,129,36.5</points>
<intersection>106 0</intersection>
<intersection>129 12</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>106,28,129,28</points>
<intersection>106 0</intersection>
<intersection>129 13</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>129,35.5,129,36.5</points>
<connection>
<GID>853</GID>
<name>ENABLE_0</name></connection>
<intersection>36.5 9</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>129,27,129,28</points>
<connection>
<GID>854</GID>
<name>ENABLE_0</name></connection>
<intersection>28 11</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>7.5,2,7.5,5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>7.5,2,28.5,2</points>
<intersection>7.5 1</intersection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,1,28.5,2</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>2 2</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>38.5,1,38.5,1</points>
<connection>
<GID>1</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-7,43,19</points>
<intersection>-7 2</intersection>
<intersection>19 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-7,43,-7</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>43,19,47,19</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-8,44,18</points>
<intersection>-8 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,18,47,18</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-8,44,-8</points>
<intersection>34 3</intersection>
<intersection>44 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-8,34,-7</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-9,45,17</points>
<intersection>-9 2</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,17,47,17</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-9,45,-9</points>
<intersection>33 3</intersection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-9,33,-7</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>-9 2</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-10,46,16</points>
<intersection>-10 2</intersection>
<intersection>16 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,-10,46,-10</points>
<intersection>32 3</intersection>
<intersection>46 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-10,32,-7</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>46,16,47,16</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-1,-18,-1,30</points>
<intersection>-18 5</intersection>
<intersection>10 45</intersection>
<intersection>14 114</intersection>
<intersection>26 44</intersection>
<intersection>30 110</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-68,-18,-1,-18</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-67 33</intersection>
<intersection>-61 123</intersection>
<intersection>-51 124</intersection>
<intersection>-41 125</intersection>
<intersection>-31 126</intersection>
<intersection>-1 3</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-67,16,-31,16</points>
<intersection>-67 33</intersection>
<intersection>-61 118</intersection>
<intersection>-51 117</intersection>
<intersection>-41 116</intersection>
<intersection>-31 115</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>-67,-18,-67,16</points>
<intersection>-18 5</intersection>
<intersection>16 20</intersection></vsegment>
<hsegment>
<ID>44</ID>
<points>-1,26,24,26</points>
<intersection>-1 3</intersection>
<intersection>8 81</intersection>
<intersection>16 85</intersection>
<intersection>24 87</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>-1,10,24.5,10</points>
<intersection>-1 3</intersection>
<intersection>8.5 89</intersection>
<intersection>16.5 93</intersection>
<intersection>24.5 95</intersection></hsegment>
<vsegment>
<ID>81</ID>
<points>8,26,8,30</points>
<connection>
<GID>116</GID>
<name>clock</name></connection>
<intersection>26 44</intersection></vsegment>
<vsegment>
<ID>85</ID>
<points>16,26,16,30</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<intersection>26 44</intersection></vsegment>
<vsegment>
<ID>87</ID>
<points>24,26,24,30</points>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<intersection>26 44</intersection></vsegment>
<vsegment>
<ID>89</ID>
<points>8.5,10,8.5,14</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>10 45</intersection></vsegment>
<vsegment>
<ID>93</ID>
<points>16.5,10,16.5,14</points>
<connection>
<GID>122</GID>
<name>clock</name></connection>
<intersection>10 45</intersection></vsegment>
<vsegment>
<ID>95</ID>
<points>24.5,10,24.5,14</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>10 45</intersection></vsegment>
<hsegment>
<ID>110</ID>
<points>-1,30,0,30</points>
<connection>
<GID>115</GID>
<name>clock</name></connection>
<intersection>-1 3</intersection></hsegment>
<hsegment>
<ID>114</ID>
<points>-1,14,0,14</points>
<connection>
<GID>120</GID>
<name>clock</name></connection>
<intersection>-1 3</intersection></hsegment>
<vsegment>
<ID>115</ID>
<points>-31,16,-31,21</points>
<intersection>16 20</intersection>
<intersection>21 120</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-41,16,-41,21</points>
<intersection>16 20</intersection>
<intersection>21 119</intersection></vsegment>
<vsegment>
<ID>117</ID>
<points>-51,16,-51,21</points>
<intersection>16 20</intersection>
<intersection>21 121</intersection></vsegment>
<vsegment>
<ID>118</ID>
<points>-61,16,-61,21</points>
<intersection>16 20</intersection>
<intersection>21 122</intersection></vsegment>
<hsegment>
<ID>119</ID>
<points>-41,21,-40,21</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>-41 116</intersection></hsegment>
<hsegment>
<ID>120</ID>
<points>-31,21,-30,21</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-31 115</intersection></hsegment>
<hsegment>
<ID>121</ID>
<points>-51,21,-50,21</points>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<intersection>-51 117</intersection></hsegment>
<hsegment>
<ID>122</ID>
<points>-61,21,-60,21</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>-61 118</intersection></hsegment>
<vsegment>
<ID>123</ID>
<points>-61,-18,-61,-13</points>
<intersection>-18 5</intersection>
<intersection>-13 127</intersection></vsegment>
<vsegment>
<ID>124</ID>
<points>-51,-18,-51,-13</points>
<intersection>-18 5</intersection>
<intersection>-13 128</intersection></vsegment>
<vsegment>
<ID>125</ID>
<points>-41,-18,-41,-13</points>
<intersection>-18 5</intersection>
<intersection>-13 129</intersection></vsegment>
<vsegment>
<ID>126</ID>
<points>-31,-18,-31,-13</points>
<intersection>-18 5</intersection>
<intersection>-13 130</intersection></vsegment>
<hsegment>
<ID>127</ID>
<points>-61,-13,-60,-13</points>
<connection>
<GID>88</GID>
<name>clock</name></connection>
<intersection>-61 123</intersection></hsegment>
<hsegment>
<ID>128</ID>
<points>-51,-13,-50,-13</points>
<connection>
<GID>94</GID>
<name>clock</name></connection>
<intersection>-51 124</intersection></hsegment>
<hsegment>
<ID>129</ID>
<points>-41,-13,-40,-13</points>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<intersection>-41 125</intersection></hsegment>
<hsegment>
<ID>130</ID>
<points>-31,-13,-30,-13</points>
<connection>
<GID>100</GID>
<name>clock</name></connection>
<intersection>-31 126</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,39,64,40.5</points>
<intersection>39 3</intersection>
<intersection>40.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,40.5,64,40.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,39,65,39</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,38,65,38</points>
<connection>
<GID>54</GID>
<name>IN_B_1</name></connection>
<intersection>63 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>63,38,63,38.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>38 1</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,36.5,64,37</points>
<intersection>36.5 2</intersection>
<intersection>37 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,36.5,64,36.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,37,65,37</points>
<connection>
<GID>54</GID>
<name>IN_B_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,34.5,64,36</points>
<intersection>34.5 2</intersection>
<intersection>36 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,34.5,64,34.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,36,65,36</points>
<connection>
<GID>54</GID>
<name>IN_B_3</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,21,64,22.5</points>
<intersection>21 3</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,22.5,64,22.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,21,65,21</points>
<connection>
<GID>39</GID>
<name>IN_B_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,20,64,20.5</points>
<intersection>20 3</intersection>
<intersection>20.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,20.5,64,20.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,20,65,20</points>
<connection>
<GID>39</GID>
<name>IN_B_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,18.5,64,19</points>
<intersection>18.5 2</intersection>
<intersection>19 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,18.5,64,18.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,19,65,19</points>
<connection>
<GID>39</GID>
<name>IN_B_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,16.5,64,18</points>
<intersection>16.5 2</intersection>
<intersection>18 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,16.5,64,16.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,18,65,18</points>
<connection>
<GID>39</GID>
<name>IN_B_3</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,3,64,4.5</points>
<intersection>3 3</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,4.5,64,4.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,3,65,3</points>
<connection>
<GID>49</GID>
<name>IN_B_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,2,64,2.5</points>
<intersection>2 3</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,2.5,64,2.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,2,65,2</points>
<connection>
<GID>49</GID>
<name>IN_B_1</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,0.5,64,1</points>
<intersection>0.5 2</intersection>
<intersection>1 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,0.5,64,0.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,1,65,1</points>
<connection>
<GID>49</GID>
<name>IN_B_2</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-1.5,64,-1.74846e-007</points>
<intersection>-1.5 2</intersection>
<intersection>-1.74846e-007 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,-1.5,64,-1.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-1.74846e-007,65,-1.74846e-007</points>
<connection>
<GID>49</GID>
<name>IN_B_3</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>56,-4,56,32</points>
<intersection>-4 9</intersection>
<intersection>14 5</intersection>
<intersection>22.5 8</intersection>
<intersection>32 10</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>56,14,65,14</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>55,22.5,56,22.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>56,-4,65,-4</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>56,32,65,32</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-5,57,31</points>
<intersection>-5 5</intersection>
<intersection>13 3</intersection>
<intersection>21.5 2</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,31,65,31</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,21.5,57,21.5</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>57,13,65,13</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>57,-5,65,-5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-6,58,30</points>
<intersection>-6 5</intersection>
<intersection>12 3</intersection>
<intersection>20.5 2</intersection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,30,65,30</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,20.5,58,20.5</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58,12,65,12</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>58,-6,65,-6</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-7,59,29</points>
<intersection>-7 5</intersection>
<intersection>11 3</intersection>
<intersection>19.5 2</intersection>
<intersection>29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,29,65,29</points>
<connection>
<GID>54</GID>
<name>IN_3</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,19.5,59,19.5</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>59,11,65,11</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>59,-7,65,-7</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,26,47,26</points>
<connection>
<GID>53</GID>
<name>IN_B_0</name></connection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,26,31,33</points>
<intersection>26 1</intersection>
<intersection>33 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>30,33,31,33</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>31 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,108.5,-10,112.5</points>
<intersection>108.5 4</intersection>
<intersection>112.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-18,112.5,-10,112.5</points>
<intersection>-18 3</intersection>
<intersection>-10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,112.5,-18,114.5</points>
<intersection>112.5 2</intersection>
<intersection>114.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11,108.5,-9,108.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-18,114.5,-17,114.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,111.5,-11,111.5</points>
<intersection>-17 3</intersection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17,109.5,-17,111.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>111.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-11,111.5,-11,115.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>111.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,106,-54,107.5</points>
<intersection>106 2</intersection>
<intersection>107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,107.5,-53,107.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,106,-54,106</points>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,105,-54,105.5</points>
<intersection>105 2</intersection>
<intersection>105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,105.5,-53,105.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,105,-54,105</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,103.5,-54,104</points>
<intersection>103.5 1</intersection>
<intersection>104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,103.5,-53,103.5</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,104,-54,104</points>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,101.5,-54,103</points>
<intersection>101.5 1</intersection>
<intersection>103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,101.5,-53,101.5</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55,103,-54,103</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,109,-29,124</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>109 6</intersection>
<intersection>113 3</intersection>
<intersection>122.5 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-29,113,-25,113</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-29,109,-25,109</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-29,122.5,-27,122.5</points>
<intersection>-29 0</intersection>
<intersection>-27 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-27,122,-27,122.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>122.5 7</intersection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,98,-60,100</points>
<connection>
<GID>129</GID>
<name>clock</name></connection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,98,-60,98</points>
<connection>
<GID>132</GID>
<name>CLK</name></connection>
<intersection>-60 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,104,-65,108</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-71,108,-65,108</points>
<intersection>-71 3</intersection>
<intersection>-65 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71,108,-71,110</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>108 2</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-72,107,-64,107</points>
<intersection>-72 3</intersection>
<intersection>-64 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-72,105,-72,107</points>
<intersection>105 17</intersection>
<intersection>107 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-64,107,-64,111</points>
<intersection>107 1</intersection>
<intersection>111 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-65,111,-59,111</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>-64 4</intersection>
<intersection>-59 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-59,109,-59,111</points>
<connection>
<GID>129</GID>
<name>count_enable</name></connection>
<intersection>111 15</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-72,105,-71,105</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-72 3</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,91,-28,111</points>
<intersection>91 4</intersection>
<intersection>98 9</intersection>
<intersection>108 2</intersection>
<intersection>111 20</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-37,108,-28,108</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>-37 3</intersection>
<intersection>-28 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-37,104,-37,108</points>
<intersection>104 24</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-78,91,-28,91</points>
<intersection>-78 18</intersection>
<intersection>-57 23</intersection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-28,98,-25,98</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-78,91,-78,111</points>
<intersection>91 4</intersection>
<intersection>111 21</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-28,111,-25,111</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-78,111,-77,111</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>-78 18</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-57,91,-57,92</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>91 4</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-43,104,-37,104</points>
<intersection>-43 25</intersection>
<intersection>-37 3</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-43,102,-43,104</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>104 24</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,100,-45,104.5</points>
<intersection>100 3</intersection>
<intersection>104.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-47,104.5,-45,104.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-45,100,-43,100</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,101,-35,105</points>
<intersection>101 4</intersection>
<intersection>105 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-44,105,-35,105</points>
<intersection>-44 3</intersection>
<intersection>-35 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-44,105,-44,107</points>
<intersection>105 2</intersection>
<intersection>107 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-37,101,-35,101</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-44,107,-43,107</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>-44 3</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-73,103,-71,103</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<connection>
<GID>139</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,112,-71,112</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,98,-58,100</points>
<connection>
<GID>129</GID>
<name>clear</name></connection>
<connection>
<GID>143</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,114,-17,114</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>-17 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-17,114,-17,116.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>114 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,107.5,-19,110</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>107.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-19,107.5,-17,107.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,95.5,-10,99.5</points>
<intersection>95.5 4</intersection>
<intersection>99.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-18,99.5,-10,99.5</points>
<intersection>-18 3</intersection>
<intersection>-10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,99.5,-18,101.5</points>
<intersection>99.5 2</intersection>
<intersection>101.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11,95.5,-9,95.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-18,101.5,-17,101.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,98.5,-11,98.5</points>
<intersection>-17 3</intersection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-17,96.5,-17,98.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>98.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-11,98.5,-11,102.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>98.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,101,-17,101</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>-17 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-17,101,-17,103.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>101 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,94.5,-19,97</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>94.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-19,94.5,-17,94.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,96,-27,118</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>96 4</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,100,-25,100</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-27,96,-25,96</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,115,-25,115</points>
<connection>
<GID>846</GID>
<name>OUT_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-79 8</intersection>
<intersection>-78 20</intersection>
<intersection>-43 62</intersection>
<intersection>-33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-33,102,-33,115</points>
<intersection>102 4</intersection>
<intersection>115 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-33,102,-25,102</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-33 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-79,90,-79,115</points>
<intersection>90 21</intersection>
<intersection>103 50</intersection>
<intersection>115 1</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>-78,113,-78,115</points>
<intersection>113 33</intersection>
<intersection>115 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-79,90,-59,90</points>
<intersection>-79 8</intersection>
<intersection>-59 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-59,90,-59,92</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>90 21</intersection></vsegment>
<hsegment>
<ID>33</ID>
<points>-78,113,-77,113</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-78 20</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>-79,103,-77,103</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-79 8</intersection></hsegment>
<vsegment>
<ID>62</ID>
<points>-43,109,-43,115</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>115 1</intersection></vsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70,80,-70,84</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-82,84,-70,84</points>
<connection>
<GID>834</GID>
<name>OUT_2</name></connection>
<intersection>-70 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>-71,78,-71,83</points>
<intersection>78 7</intersection>
<intersection>83 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-71,78,-70,78</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>-71 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-82,83,-71,83</points>
<connection>
<GID>834</GID>
<name>OUT_1</name></connection>
<intersection>-71 6</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64,79,-62,79</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<connection>
<GID>407</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,78,-55,83</points>
<intersection>78 2</intersection>
<intersection>83 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-56,78,-55,78</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55,83,-54,83</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-82,82,-72,82</points>
<connection>
<GID>834</GID>
<name>OUT_0</name></connection>
<intersection>-72 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-72,71,-72,82</points>
<intersection>71 10</intersection>
<intersection>82 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-72,71,-70,71</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>-72 9</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,71,-63,77</points>
<intersection>71 2</intersection>
<intersection>77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,77,-62,77</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64,71,-63,71</points>
<connection>
<GID>415</GID>
<name>OUT_0</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,80,-40,83</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,80,-40,80</points>
<intersection>-46 3</intersection>
<intersection>-40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-46,77,-46,80</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>80 1</intersection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-48,84,-46,84</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<connection>
<GID>410</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-48,64,-46,64</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-72,62,-46,62</points>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<intersection>-59 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-59,62,-59,75</points>
<intersection>62 1</intersection>
<intersection>75 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-59,75,-46,75</points>
<connection>
<GID>417</GID>
<name>IN_1</name></connection>
<intersection>-59 3</intersection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,79,-47,82</points>
<intersection>79 2</intersection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,82,-46,82</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>-47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,79,-39,79</points>
<intersection>-47 0</intersection>
<intersection>-39 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-39,76,-39,79</points>
<intersection>76 4</intersection>
<intersection>79 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-40,76,-35,76</points>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<connection>
<GID>417</GID>
<name>OUT</name></connection>
<intersection>-39 3</intersection>
<intersection>-38 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-38,70,-38,76</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>76 4</intersection></vsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,68,-38,68</points>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection>
<connection>
<GID>429</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32,69,-30,69</points>
<connection>
<GID>429</GID>
<name>OUT</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,60,-35,63</points>
<intersection>60 1</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,60,-30,60</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-40,63,-35,63</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,61,-23,64</points>
<intersection>61 2</intersection>
<intersection>64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31,64,-23,64</points>
<intersection>-31 3</intersection>
<intersection>-23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24,61,-21,61</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<connection>
<GID>422</GID>
<name>N_in0</name></connection>
<intersection>-23 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-31,64,-31,67</points>
<intersection>64 1</intersection>
<intersection>67 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-31,67,-30,67</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<intersection>-31 3</intersection></hsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,85,-54,85</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<connection>
<GID>834</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,65,-24,68</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,65,-24,65</points>
<intersection>-30 3</intersection>
<intersection>-24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30,62,-30,65</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>65 1</intersection></vsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>232.5,58.5,232.5,58.5</points>
<connection>
<GID>542</GID>
<name>clock</name></connection>
<connection>
<GID>543</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>232.5,69.5,232.5,69.5</points>
<connection>
<GID>542</GID>
<name>load</name></connection>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,50,221.5,67.5</points>
<intersection>50 2</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221.5,67.5,229.5,67.5</points>
<connection>
<GID>542</GID>
<name>IN_7</name></connection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,50,221.5,50</points>
<connection>
<GID>506</GID>
<name>OUT</name></connection>
<intersection>221.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,54,222.5,66.5</points>
<intersection>54 2</intersection>
<intersection>66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,66.5,229.5,66.5</points>
<connection>
<GID>542</GID>
<name>IN_6</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,54,222.5,54</points>
<connection>
<GID>505</GID>
<name>OUT</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,58,223.5,65.5</points>
<intersection>58 2</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,65.5,229.5,65.5</points>
<connection>
<GID>542</GID>
<name>IN_5</name></connection>
<intersection>223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,58,223.5,58</points>
<connection>
<GID>504</GID>
<name>OUT</name></connection>
<intersection>223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>224.5,64.5,229.5,64.5</points>
<connection>
<GID>542</GID>
<name>IN_4</name></connection>
<intersection>224.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>224.5,62,224.5,64.5</points>
<intersection>62 4</intersection>
<intersection>64.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>220.5,62,224.5,62</points>
<connection>
<GID>503</GID>
<name>OUT</name></connection>
<intersection>224.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225.5,63.5,229.5,63.5</points>
<connection>
<GID>542</GID>
<name>IN_3</name></connection>
<intersection>225.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>225.5,63.5,225.5,66</points>
<intersection>63.5 1</intersection>
<intersection>66 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>220.5,66,225.5,66</points>
<connection>
<GID>502</GID>
<name>OUT</name></connection>
<intersection>225.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,62.5,226.5,70</points>
<intersection>62.5 1</intersection>
<intersection>70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,62.5,229.5,62.5</points>
<connection>
<GID>542</GID>
<name>IN_2</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,70,226.5,70</points>
<connection>
<GID>501</GID>
<name>OUT</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>175,123.5,175,129</points>
<intersection>123.5 34</intersection>
<intersection>129 16</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>131.5,129,176.5,129</points>
<intersection>131.5 59</intersection>
<intersection>175 5</intersection>
<intersection>176.5 58</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>175,123.5,175.5,123.5</points>
<intersection>175 5</intersection>
<intersection>175.5 41</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>175.5,122,175.5,123.5</points>
<connection>
<GID>444</GID>
<name>load</name></connection>
<intersection>123.5 34</intersection></vsegment>
<vsegment>
<ID>58</ID>
<points>176.5,126,176.5,129</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>129 16</intersection></vsegment>
<vsegment>
<ID>59</ID>
<points>131.5,125,131.5,129</points>
<connection>
<GID>857</GID>
<name>OUT_0</name></connection>
<intersection>129 16</intersection></vsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,122,176.5,122</points>
<connection>
<GID>441</GID>
<name>OUT_0</name></connection>
<connection>
<GID>444</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,122,177.5,131</points>
<connection>
<GID>444</GID>
<name>count_up</name></connection>
<intersection>131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,131,177.5,131</points>
<connection>
<GID>856</GID>
<name>OUT_0</name></connection>
<intersection>140.5 2</intersection>
<intersection>177.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>140.5,131,140.5,149</points>
<intersection>131 1</intersection>
<intersection>137 6</intersection>
<intersection>149 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>140.5,137,144.5,137</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>140.5 2</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>140.5,149,150.5,149</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>140.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,82,189.5,150</points>
<intersection>82 3</intersection>
<intersection>120 2</intersection>
<intersection>150 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,150,190.5,150</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180.5,120,189.5,120</points>
<connection>
<GID>444</GID>
<name>OUT_7</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>189.5,82,194.5,82</points>
<connection>
<GID>540</GID>
<name>IN_1</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,86,188.5,154</points>
<intersection>86 3</intersection>
<intersection>119 2</intersection>
<intersection>154 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,154,190.5,154</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180.5,119,188.5,119</points>
<connection>
<GID>444</GID>
<name>OUT_6</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>188.5,86,194.5,86</points>
<connection>
<GID>539</GID>
<name>IN_1</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,90,187.5,158</points>
<intersection>90 4</intersection>
<intersection>118 2</intersection>
<intersection>158 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187.5,158,190.5,158</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180.5,118,187.5,118</points>
<connection>
<GID>444</GID>
<name>OUT_5</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>187.5,90,194.5,90</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,94,186.5,162</points>
<intersection>94 4</intersection>
<intersection>117 2</intersection>
<intersection>162 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,162,190.5,162</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180.5,117,186.5,117</points>
<connection>
<GID>444</GID>
<name>OUT_4</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>186.5,94,194.5,94</points>
<connection>
<GID>537</GID>
<name>IN_1</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,98,185.5,166</points>
<intersection>98 4</intersection>
<intersection>116 1</intersection>
<intersection>166 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,116,185.5,116</points>
<connection>
<GID>444</GID>
<name>OUT_3</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185.5,166,190.5,166</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185.5,98,194.5,98</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,102,184.5,170</points>
<intersection>102 3</intersection>
<intersection>115 1</intersection>
<intersection>170 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,115,184.5,115</points>
<connection>
<GID>444</GID>
<name>OUT_2</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,170,190.5,170</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>184.5,102,194.5,102</points>
<connection>
<GID>535</GID>
<name>IN_1</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,106,183.5,174</points>
<intersection>106 3</intersection>
<intersection>114 1</intersection>
<intersection>174 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,114,183.5,114</points>
<connection>
<GID>444</GID>
<name>OUT_1</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,174,190.5,174</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>183.5,106,194.5,106</points>
<connection>
<GID>534</GID>
<name>IN_1</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182.5,110,182.5,178</points>
<intersection>110 3</intersection>
<intersection>113 1</intersection>
<intersection>178 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,113,182.5,113</points>
<connection>
<GID>444</GID>
<name>OUT_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182.5,178,190.5,178</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<intersection>182.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>182.5,110,194.5,110</points>
<connection>
<GID>533</GID>
<name>IN_1</name></connection>
<intersection>182.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,61.5,227.5,74</points>
<intersection>61.5 1</intersection>
<intersection>74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,61.5,229.5,61.5</points>
<connection>
<GID>542</GID>
<name>IN_1</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,74,227.5,74</points>
<connection>
<GID>500</GID>
<name>OUT</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,60.5,228.5,78</points>
<intersection>60.5 3</intersection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>220.5,78,228.5,78</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>228.5,60.5,229.5,60.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>255.5,120.5,255.5,120.5</points>
<connection>
<GID>546</GID>
<name>load</name></connection>
<connection>
<GID>548</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>255.5,109.5,255.5,109.5</points>
<connection>
<GID>546</GID>
<name>clock</name></connection>
<connection>
<GID>547</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,101,244.5,118.5</points>
<intersection>101 2</intersection>
<intersection>118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,118.5,252.5,118.5</points>
<connection>
<GID>546</GID>
<name>IN_7</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,101,244.5,101</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,105,245.5,117.5</points>
<intersection>105 2</intersection>
<intersection>117.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,117.5,252.5,117.5</points>
<connection>
<GID>546</GID>
<name>IN_6</name></connection>
<intersection>245.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,105,245.5,105</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,109,246.5,116.5</points>
<intersection>109 2</intersection>
<intersection>116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246.5,116.5,252.5,116.5</points>
<connection>
<GID>546</GID>
<name>IN_5</name></connection>
<intersection>246.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,109,246.5,109</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>246.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247.5,113,247.5,115.5</points>
<intersection>113 2</intersection>
<intersection>115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247.5,115.5,252.5,115.5</points>
<connection>
<GID>546</GID>
<name>IN_4</name></connection>
<intersection>247.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,113,247.5,113</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>247.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248.5,114.5,248.5,117</points>
<intersection>114.5 3</intersection>
<intersection>117 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>243.5,117,248.5,117</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>248.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>248.5,114.5,252.5,114.5</points>
<connection>
<GID>546</GID>
<name>IN_3</name></connection>
<intersection>248.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,113.5,249.5,121</points>
<intersection>113.5 1</intersection>
<intersection>121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249.5,113.5,252.5,113.5</points>
<connection>
<GID>546</GID>
<name>IN_2</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,121,249.5,121</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250.5,112.5,250.5,125</points>
<intersection>112.5 1</intersection>
<intersection>125 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250.5,112.5,252.5,112.5</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<intersection>250.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,125,250.5,125</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>250.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251.5,111.5,251.5,129</points>
<intersection>111.5 1</intersection>
<intersection>129 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251.5,111.5,252.5,111.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>251.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,129,251.5,129</points>
<connection>
<GID>458</GID>
<name>OUT</name></connection>
<intersection>251.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,171.5,232.5,171.5</points>
<connection>
<GID>541</GID>
<name>load</name></connection>
<connection>
<GID>545</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,160.5,232.5,160.5</points>
<connection>
<GID>541</GID>
<name>clock</name></connection>
<connection>
<GID>544</GID>
<name>CLK</name></connection></vsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,152,228.5,169.5</points>
<intersection>152 2</intersection>
<intersection>169.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,169.5,229.5,169.5</points>
<connection>
<GID>541</GID>
<name>IN_7</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,152,228.5,152</points>
<connection>
<GID>474</GID>
<name>OUT</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,156,227.5,168.5</points>
<intersection>156 2</intersection>
<intersection>168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,168.5,229.5,168.5</points>
<connection>
<GID>541</GID>
<name>IN_6</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,156,227.5,156</points>
<connection>
<GID>473</GID>
<name>OUT</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,160,226.5,167.5</points>
<intersection>160 2</intersection>
<intersection>167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,167.5,229.5,167.5</points>
<connection>
<GID>541</GID>
<name>IN_5</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,160,226.5,160</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,164,225.5,166.5</points>
<intersection>164 2</intersection>
<intersection>166.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,166.5,229.5,166.5</points>
<connection>
<GID>541</GID>
<name>IN_4</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,164,225.5,164</points>
<connection>
<GID>471</GID>
<name>OUT</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,165.5,224.5,168</points>
<intersection>165.5 1</intersection>
<intersection>168 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224.5,165.5,229.5,165.5</points>
<connection>
<GID>541</GID>
<name>IN_3</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,168,224.5,168</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<intersection>224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,164.5,223.5,172</points>
<intersection>164.5 1</intersection>
<intersection>172 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,164.5,229.5,164.5</points>
<connection>
<GID>541</GID>
<name>IN_2</name></connection>
<intersection>223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,172,223.5,172</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<intersection>223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,163.5,222.5,176</points>
<intersection>163.5 1</intersection>
<intersection>176 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,163.5,229.5,163.5</points>
<connection>
<GID>541</GID>
<name>IN_1</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,176,222.5,176</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,162.5,221.5,180</points>
<intersection>162.5 1</intersection>
<intersection>180 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221.5,162.5,229.5,162.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,180,221.5,180</points>
<connection>
<GID>466</GID>
<name>OUT</name></connection>
<intersection>221.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236.5,84,236.5,100</points>
<intersection>84 2</intersection>
<intersection>100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,100,237.5,100</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>236.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,84,236.5,84</points>
<connection>
<GID>498</GID>
<name>OUT</name></connection>
<intersection>236.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,88,235.5,104</points>
<intersection>88 2</intersection>
<intersection>104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235.5,104,237.5,104</points>
<connection>
<GID>464</GID>
<name>IN_1</name></connection>
<intersection>235.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,88,235.5,88</points>
<connection>
<GID>497</GID>
<name>OUT</name></connection>
<intersection>235.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,92,234.5,108</points>
<intersection>92 2</intersection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,108,237.5,108</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,92,234.5,92</points>
<connection>
<GID>496</GID>
<name>OUT</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233.5,96,233.5,112</points>
<intersection>96 2</intersection>
<intersection>112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>233.5,112,237.5,112</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<intersection>233.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,96,233.5,96</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<intersection>233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,100,232.5,116</points>
<intersection>100 2</intersection>
<intersection>116 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>232.5,116,237.5,116</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,100,232.5,100</points>
<connection>
<GID>494</GID>
<name>OUT</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,104,231.5,120</points>
<intersection>104 2</intersection>
<intersection>120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,120,237.5,120</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>231.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,104,231.5,104</points>
<connection>
<GID>493</GID>
<name>OUT</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,108,230.5,124</points>
<intersection>108 2</intersection>
<intersection>124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,124,237.5,124</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<intersection>230.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,108,230.5,108</points>
<connection>
<GID>492</GID>
<name>OUT</name></connection>
<intersection>230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,112,229.5,128</points>
<intersection>112 2</intersection>
<intersection>128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,128,237.5,128</points>
<connection>
<GID>458</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,112,229.5,112</points>
<connection>
<GID>490</GID>
<name>OUT</name></connection>
<intersection>229.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,130,228.5,146</points>
<intersection>130 1</intersection>
<intersection>146 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>228.5,130,237.5,130</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>228.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,146,228.5,146</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<intersection>228.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227.5,126,227.5,142</points>
<intersection>126 1</intersection>
<intersection>142 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227.5,126,237.5,126</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>227.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>220.5,142,227.5,142</points>
<connection>
<GID>476</GID>
<name>OUT</name></connection>
<intersection>227.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,141,139.5,145</points>
<intersection>141 4</intersection>
<intersection>143 5</intersection>
<intersection>145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,145,142.5,145</points>
<connection>
<GID>447</GID>
<name>J</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>139.5,141,142.5,141</points>
<connection>
<GID>447</GID>
<name>K</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>138.5,143,139.5,143</points>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,135,178.5,135</points>
<intersection>141.5 27</intersection>
<intersection>166.5 28</intersection>
<intersection>178.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>178.5,122,178.5,135</points>
<connection>
<GID>444</GID>
<name>carry_out</name></connection>
<intersection>135 1</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>141.5,135,141.5,143</points>
<intersection>135 1</intersection>
<intersection>143 29</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>166.5,135,166.5,143</points>
<intersection>135 1</intersection>
<intersection>143 30</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>141.5,143,142.5,143</points>
<connection>
<GID>447</GID>
<name>clock</name></connection>
<intersection>141.5 27</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>166.5,143,167.5,143</points>
<connection>
<GID>448</GID>
<name>clock</name></connection>
<intersection>166.5 28</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148.5,137,150.5,137</points>
<connection>
<GID>453</GID>
<name>OUT_0</name></connection>
<connection>
<GID>452</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,122,226.5,138</points>
<intersection>122 1</intersection>
<intersection>138 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226.5,122,237.5,122</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,138,226.5,138</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<intersection>226.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,139,149.5,141</points>
<intersection>139 6</intersection>
<intersection>141 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148.5,141,149.5,141</points>
<connection>
<GID>447</GID>
<name>nQ</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>149.5,139,150.5,139</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,118,225.5,134</points>
<intersection>118 1</intersection>
<intersection>134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,118,237.5,118</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,134,225.5,134</points>
<connection>
<GID>478</GID>
<name>OUT</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,144,157.5,148</points>
<intersection>144 10</intersection>
<intersection>148 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>156.5,148,157.5,148</points>
<connection>
<GID>451</GID>
<name>OUT</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>157.5,144,158.5,144</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>157.5,138,157.5,142</points>
<intersection>138 15</intersection>
<intersection>142 16</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>156.5,138,157.5,138</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>157.5 5</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>157.5,142,158.5,142</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<intersection>157.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>165.5,141,165.5,145</points>
<intersection>141 10</intersection>
<intersection>143 15</intersection>
<intersection>145 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>165.5,145,167.5,145</points>
<connection>
<GID>448</GID>
<name>J</name></connection>
<intersection>165.5 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>165.5,141,167.5,141</points>
<connection>
<GID>448</GID>
<name>K</name></connection>
<intersection>165.5 7</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>164.5,143,165.5,143</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<intersection>165.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224.5,114,224.5,130</points>
<intersection>114 3</intersection>
<intersection>130 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>220.5,130,224.5,130</points>
<connection>
<GID>479</GID>
<name>OUT</name></connection>
<intersection>224.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>224.5,114,237.5,114</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,110,223.5,126</points>
<intersection>110 1</intersection>
<intersection>126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>223.5,110,237.5,110</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>223.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,126,223.5,126</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<intersection>223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,106,222.5,122</points>
<intersection>106 1</intersection>
<intersection>122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,106,237.5,106</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,122,222.5,122</points>
<connection>
<GID>481</GID>
<name>OUT</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,102,221.5,118</points>
<intersection>102 1</intersection>
<intersection>118 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>221.5,102,237.5,102</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,118,221.5,118</points>
<connection>
<GID>482</GID>
<name>OUT</name></connection>
<intersection>221.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,110,177.5,111</points>
<connection>
<GID>432</GID>
<name>OUT_0</name></connection>
<connection>
<GID>444</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,181,214.5,181</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<connection>
<GID>467</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>209.5,145,209.5,179</points>
<intersection>145 19</intersection>
<intersection>179 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>200.5,179,214.5,179</points>
<connection>
<GID>523</GID>
<name>OUT</name></connection>
<connection>
<GID>466</GID>
<name>IN_1</name></connection>
<intersection>209.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>209.5,145,214.5,145</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>209.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,141,208.5,175</points>
<intersection>141 3</intersection>
<intersection>175 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,175,214.5,175</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>208.5,141,214.5,141</points>
<connection>
<GID>476</GID>
<name>IN_1</name></connection>
<intersection>208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,137,207.5,171</points>
<intersection>137 3</intersection>
<intersection>171 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,171,214.5,171</points>
<connection>
<GID>525</GID>
<name>OUT</name></connection>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,137,214.5,137</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>206.5,133,206.5,167</points>
<intersection>133 5</intersection>
<intersection>167 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>206.5,133,214.5,133</points>
<connection>
<GID>478</GID>
<name>IN_1</name></connection>
<intersection>206.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,167,214.5,167</points>
<connection>
<GID>526</GID>
<name>OUT</name></connection>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>206.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>205.5,129,205.5,163</points>
<intersection>129 4</intersection>
<intersection>163 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>205.5,129,214.5,129</points>
<connection>
<GID>479</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,163,214.5,163</points>
<connection>
<GID>527</GID>
<name>OUT</name></connection>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,159,214.5,159</points>
<connection>
<GID>528</GID>
<name>OUT</name></connection>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>205.5,125,205.5,159</points>
<intersection>125 4</intersection>
<intersection>159 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>205.5,125,214.5,125</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,155,214.5,155</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>473</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>204.5,121,204.5,155</points>
<intersection>121 4</intersection>
<intersection>155 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>204.5,121,214.5,121</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>202.5,117,202.5,151</points>
<intersection>117 4</intersection>
<intersection>151 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>202.5,117,214.5,117</points>
<connection>
<GID>482</GID>
<name>IN_1</name></connection>
<intersection>202.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>200.5,151,214.5,151</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>202.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,153,214.5,153</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<connection>
<GID>489</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,157,214.5,157</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>488</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,161,214.5,161</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<connection>
<GID>487</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,165,214.5,165</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,169,214.5,169</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<connection>
<GID>485</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,173,214.5,173</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<connection>
<GID>484</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,177,214.5,177</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<connection>
<GID>483</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,113,214.5,113</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<connection>
<GID>491</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>508</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>209.5,77,209.5,111</points>
<intersection>77 19</intersection>
<intersection>111 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>200.5,111,214.5,111</points>
<connection>
<GID>533</GID>
<name>OUT</name></connection>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<intersection>209.5 3</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>209.5,77,214.5,77</points>
<connection>
<GID>499</GID>
<name>IN_1</name></connection>
<intersection>209.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208.5,73,208.5,107</points>
<intersection>73 3</intersection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,107,214.5,107</points>
<connection>
<GID>534</GID>
<name>OUT</name></connection>
<connection>
<GID>492</GID>
<name>IN_1</name></connection>
<intersection>208.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>208.5,73,214.5,73</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>208.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,69,207.5,103</points>
<intersection>69 3</intersection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,103,214.5,103</points>
<connection>
<GID>535</GID>
<name>OUT</name></connection>
<connection>
<GID>493</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207.5,69,214.5,69</points>
<connection>
<GID>501</GID>
<name>IN_1</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>206.5,65,206.5,99</points>
<intersection>65 5</intersection>
<intersection>99 8</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>206.5,65,214.5,65</points>
<connection>
<GID>502</GID>
<name>IN_1</name></connection>
<intersection>206.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,99,214.5,99</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>206.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>205.5,61,205.5,95</points>
<intersection>61 4</intersection>
<intersection>95 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>205.5,61,214.5,61</points>
<connection>
<GID>503</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,95,214.5,95</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<connection>
<GID>495</GID>
<name>IN_1</name></connection>
<intersection>205.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>204.5,57,204.5,91</points>
<intersection>57 4</intersection>
<intersection>91 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>204.5,57,214.5,57</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,91,214.5,91</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<connection>
<GID>496</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,87,214.5,87</points>
<connection>
<GID>539</GID>
<name>OUT</name></connection>
<connection>
<GID>497</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>204.5,53,204.5,87</points>
<intersection>53 4</intersection>
<intersection>87 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>204.5,53,214.5,53</points>
<connection>
<GID>505</GID>
<name>IN_1</name></connection>
<intersection>204.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>202.5,49,202.5,83</points>
<intersection>49 4</intersection>
<intersection>83 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>202.5,49,214.5,49</points>
<connection>
<GID>506</GID>
<name>IN_1</name></connection>
<intersection>202.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>200.5,83,214.5,83</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<connection>
<GID>498</GID>
<name>IN_1</name></connection>
<intersection>202.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,85,214.5,85</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<connection>
<GID>513</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,51,201.5,185.5</points>
<intersection>51 18</intersection>
<intersection>55 17</intersection>
<intersection>59 16</intersection>
<intersection>63 15</intersection>
<intersection>67 14</intersection>
<intersection>71 13</intersection>
<intersection>75 12</intersection>
<intersection>79 11</intersection>
<intersection>85 2</intersection>
<intersection>89 9</intersection>
<intersection>93 8</intersection>
<intersection>97 7</intersection>
<intersection>101 6</intersection>
<intersection>105 5</intersection>
<intersection>109 4</intersection>
<intersection>113 3</intersection>
<intersection>119 38</intersection>
<intersection>123 37</intersection>
<intersection>127 36</intersection>
<intersection>131 35</intersection>
<intersection>135 34</intersection>
<intersection>139 33</intersection>
<intersection>143 32</intersection>
<intersection>147 31</intersection>
<intersection>153 22</intersection>
<intersection>157 29</intersection>
<intersection>161 28</intersection>
<intersection>165 27</intersection>
<intersection>169 26</intersection>
<intersection>173 25</intersection>
<intersection>177 24</intersection>
<intersection>181 23</intersection>
<intersection>185.5 48</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>201.5,85,210.5,85</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>201.5,113,210.5,113</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>201.5,109,210.5,109</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>201.5,105,210.5,105</points>
<connection>
<GID>508</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>201.5,101,210.5,101</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>201.5,97,210.5,97</points>
<connection>
<GID>510</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>201.5,93,210.5,93</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>201.5,89,210.5,89</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>201.5,79,214.5,79</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>201.5,75,214.5,75</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>201.5,71,214.5,71</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>201.5,67,214.5,67</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>201.5,63,214.5,63</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>201.5,59,214.5,59</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>201.5,55,214.5,55</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>201.5,51,214.5,51</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>201.5,153,210.5,153</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>201.5,181,210.5,181</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>201.5,177,210.5,177</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>201.5,173,210.5,173</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>201.5,169,210.5,169</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>201.5,165,210.5,165</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>201.5,161,210.5,161</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>201.5,157,210.5,157</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>201.5,147,214.5,147</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>201.5,143,214.5,143</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>201.5,139,214.5,139</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>201.5,135,214.5,135</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>201.5,131,214.5,131</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>201.5,127,214.5,127</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>201.5,123,214.5,123</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>38</ID>
<points>201.5,119,214.5,119</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>201.5 0</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>174.5,185.5,201.5,185.5</points>
<intersection>174.5 49</intersection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>49</ID>
<points>174.5,145,174.5,185.5</points>
<intersection>145 52</intersection>
<intersection>185.5 48</intersection></vsegment>
<hsegment>
<ID>52</ID>
<points>173.5,145,174.5,145</points>
<connection>
<GID>448</GID>
<name>Q</name></connection>
<intersection>174.5 49</intersection></hsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,89,214.5,89</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<connection>
<GID>512</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,93,214.5,93</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<connection>
<GID>511</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,97,214.5,97</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<connection>
<GID>510</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,101,214.5,101</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,105,214.5,105</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<connection>
<GID>508</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,109,214.5,109</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<connection>
<GID>507</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,178,194.5,178</points>
<connection>
<GID>515</GID>
<name>OUT_0</name></connection>
<connection>
<GID>523</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,174,194.5,174</points>
<connection>
<GID>516</GID>
<name>OUT_0</name></connection>
<connection>
<GID>524</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,170,194.5,170</points>
<connection>
<GID>517</GID>
<name>OUT_0</name></connection>
<connection>
<GID>525</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,166,194.5,166</points>
<connection>
<GID>518</GID>
<name>OUT_0</name></connection>
<connection>
<GID>526</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,162,194.5,162</points>
<connection>
<GID>519</GID>
<name>OUT_0</name></connection>
<connection>
<GID>527</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,158,194.5,158</points>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection>
<connection>
<GID>528</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,154,194.5,154</points>
<connection>
<GID>521</GID>
<name>OUT_0</name></connection>
<connection>
<GID>529</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,150,194.5,150</points>
<connection>
<GID>522</GID>
<name>OUT_0</name></connection>
<connection>
<GID>530</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180.5,180,194.5,180</points>
<connection>
<GID>531</GID>
<name>OUT_0</name></connection>
<connection>
<GID>523</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>182.5,152,182.5,180</points>
<intersection>152 4</intersection>
<intersection>156 10</intersection>
<intersection>160 9</intersection>
<intersection>164 8</intersection>
<intersection>168 7</intersection>
<intersection>172 6</intersection>
<intersection>176 5</intersection>
<intersection>180 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>182.5,152,194.5,152</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>182.5,176,194.5,176</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>182.5,172,194.5,172</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>182.5,168,194.5,168</points>
<connection>
<GID>526</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>182.5,164,194.5,164</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>182.5,160,194.5,160</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>182.5,156,194.5,156</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>182.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149.5,151,181.5,151</points>
<intersection>149.5 45</intersection>
<intersection>175.5 12</intersection>
<intersection>181.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>181.5,84,181.5,151</points>
<intersection>84 4</intersection>
<intersection>88 10</intersection>
<intersection>92 9</intersection>
<intersection>96 8</intersection>
<intersection>100 7</intersection>
<intersection>104 6</intersection>
<intersection>108 5</intersection>
<intersection>112 28</intersection>
<intersection>151 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>181.5,84,194.5,84</points>
<connection>
<GID>540</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>181.5,108,194.5,108</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>181.5,104,194.5,104</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>181.5,100,194.5,100</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>181.5,96,194.5,96</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>181.5,92,194.5,92</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>181.5,88,194.5,88</points>
<connection>
<GID>539</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>175.5,151,175.5,180</points>
<intersection>151 1</intersection>
<intersection>180 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>175.5,180,176.5,180</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>175.5 12</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>181.5,112,194.5,112</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>181.5 3</intersection></hsegment>
<vsegment>
<ID>45</ID>
<points>149.5,145,149.5,151</points>
<intersection>145 47</intersection>
<intersection>147 48</intersection>
<intersection>151 1</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>148.5,145,149.5,145</points>
<connection>
<GID>447</GID>
<name>Q</name></connection>
<intersection>149.5 45</intersection></hsegment>
<hsegment>
<ID>48</ID>
<points>149.5,147,150.5,147</points>
<connection>
<GID>451</GID>
<name>IN_1</name></connection>
<intersection>149.5 45</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>250.5,27,278.5,27</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>250.5 29</intersection>
<intersection>258 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>258,-29,258,27</points>
<intersection>-29 15</intersection>
<intersection>-21 17</intersection>
<intersection>-13 18</intersection>
<intersection>-5 19</intersection>
<intersection>3 20</intersection>
<intersection>11 21</intersection>
<intersection>19 16</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>258,-29,278.5,-29</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>258,19,278.5,19</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>258,-21,278.5,-21</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>258,-13,278.5,-13</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>258,-5,278.5,-5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>258,3,278.5,3</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>258,11,278.5,11</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>258 13</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>250.5,-11,250.5,27</points>
<intersection>-11 30</intersection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>248,-11,250.5,-11</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<intersection>250.5 29</intersection></hsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>184,-3,185,-3</points>
<connection>
<GID>581</GID>
<name>IN_1</name></connection>
<connection>
<GID>578</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>187,-3,188,-3</points>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<connection>
<GID>580</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>19</ID>
<points>253,-27,253,31.5</points>
<intersection>-27 79</intersection>
<intersection>31.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>253,31.5,369.5,31.5</points>
<intersection>253 19</intersection>
<intersection>369.5 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>369.5,-68.5,369.5,31.5</points>
<intersection>-68.5 47</intersection>
<intersection>-8.5 69</intersection>
<intersection>31.5 24</intersection></vsegment>
<hsegment>
<ID>47</ID>
<points>369.5,-68.5,439,-68.5</points>
<intersection>369.5 36</intersection>
<intersection>384.5 77</intersection>
<intersection>393.5 59</intersection>
<intersection>402.5 60</intersection>
<intersection>412 61</intersection>
<intersection>421 63</intersection>
<intersection>430 64</intersection>
<intersection>439 65</intersection></hsegment>
<vsegment>
<ID>59</ID>
<points>393.5,-69,393.5,-68.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<vsegment>
<ID>60</ID>
<points>402.5,-69,402.5,-68.5</points>
<connection>
<GID>677</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>412,-69,412,-68.5</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<vsegment>
<ID>63</ID>
<points>421,-69,421,-68.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<vsegment>
<ID>64</ID>
<points>430,-69,430,-68.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<vsegment>
<ID>65</ID>
<points>439,-69,439,-68.5</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<hsegment>
<ID>69</ID>
<points>369.5,-8.5,437.5,-8.5</points>
<intersection>369.5 36</intersection>
<intersection>383 76</intersection>
<intersection>392 75</intersection>
<intersection>401 74</intersection>
<intersection>410.5 73</intersection>
<intersection>419.5 72</intersection>
<intersection>428.5 71</intersection>
<intersection>437.5 70</intersection></hsegment>
<vsegment>
<ID>70</ID>
<points>437.5,-9.5,437.5,-8.5</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>71</ID>
<points>428.5,-9.5,428.5,-8.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>72</ID>
<points>419.5,-9.5,419.5,-8.5</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>73</ID>
<points>410.5,-9.5,410.5,-8.5</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>74</ID>
<points>401,-9.5,401,-8.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>75</ID>
<points>392,-9.5,392,-8.5</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>76</ID>
<points>383,-9.5,383,-8.5</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>-8.5 69</intersection></vsegment>
<vsegment>
<ID>77</ID>
<points>384.5,-69,384.5,-68.5</points>
<connection>
<GID>667</GID>
<name>IN_0</name></connection>
<intersection>-68.5 47</intersection></vsegment>
<hsegment>
<ID>79</ID>
<points>206,-27,253,-27</points>
<connection>
<GID>659</GID>
<name>OUT_0</name></connection>
<intersection>253 19</intersection></hsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-8.5,181.5,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-8.5,184.5,-8.5</points>
<intersection>181.5 0</intersection>
<intersection>184.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,3,183,3</points>
<connection>
<GID>578</GID>
<name>IN_1</name></connection>
<intersection>181.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>184.5,-11,184.5,-8.5</points>
<connection>
<GID>577</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>193,-3,194,-3</points>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<connection>
<GID>587</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>196,-3,197,-3</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<connection>
<GID>588</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-8.5,190.5,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190.5,-8.5,193.5,-8.5</points>
<intersection>190.5 0</intersection>
<intersection>193.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190.5,3,192,3</points>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<intersection>190.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>193.5,-11,193.5,-8.5</points>
<connection>
<GID>585</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>202,-3,203,-3</points>
<connection>
<GID>593</GID>
<name>IN_1</name></connection>
<connection>
<GID>591</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>205,-3,206,-3</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<connection>
<GID>592</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199.5,-8.5,199.5,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199.5,-8.5,202.5,-8.5</points>
<intersection>199.5 0</intersection>
<intersection>202.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,3,201,3</points>
<connection>
<GID>591</GID>
<name>IN_1</name></connection>
<intersection>199.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>202.5,-11,202.5,-8.5</points>
<connection>
<GID>590</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>211.5,-3,212.5,-3</points>
<connection>
<GID>597</GID>
<name>IN_1</name></connection>
<connection>
<GID>595</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>214.5,-3,215.5,-3</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<connection>
<GID>596</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-8.5,209,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,-8.5,212,-8.5</points>
<intersection>209 0</intersection>
<intersection>212 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,3,210.5,3</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<intersection>209 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>212,-11,212,-8.5</points>
<connection>
<GID>594</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>220.5,-3,221.5,-3</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<connection>
<GID>599</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>223.5,-3,224.5,-3</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<connection>
<GID>600</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-8.5,218,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-8.5,221,-8.5</points>
<intersection>218 0</intersection>
<intersection>221 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>218,3,219.5,3</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>218 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>221,-11,221,-8.5</points>
<connection>
<GID>598</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>229.5,-3,230.5,-3</points>
<connection>
<GID>605</GID>
<name>IN_1</name></connection>
<connection>
<GID>603</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>561</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>232.5,-3,233.5,-3</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<connection>
<GID>604</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-8.5,227,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>227,-8.5,230,-8.5</points>
<intersection>227 0</intersection>
<intersection>230 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>227,3,228.5,3</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<intersection>227 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>230,-11,230,-8.5</points>
<connection>
<GID>602</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>238.5,-3,239.5,-3</points>
<connection>
<GID>609</GID>
<name>IN_1</name></connection>
<connection>
<GID>607</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>241.5,-3,242.5,-3</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<connection>
<GID>608</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>236,-8.5,236,3</points>
<intersection>-8.5 1</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236,-8.5,239,-8.5</points>
<intersection>236 0</intersection>
<intersection>239 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>236,3,237.5,3</points>
<connection>
<GID>607</GID>
<name>IN_1</name></connection>
<intersection>236 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239,-11,239,-8.5</points>
<connection>
<GID>606</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-11,176,6.5</points>
<intersection>-11 4</intersection>
<intersection>6.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>172.5,6.5,176,6.5</points>
<connection>
<GID>613</GID>
<name>OUT_0</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>176,-11,178.5,-11</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,3,187,7.5</points>
<connection>
<GID>580</GID>
<name>IN_1</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,7.5,187,7.5</points>
<connection>
<GID>613</GID>
<name>OUT_1</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-11,186,-9</points>
<connection>
<GID>581</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,-11,187.5,-11</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204,-11,204,-9</points>
<connection>
<GID>593</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204,-11,206,-11</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<intersection>204 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195,-11,195,-9</points>
<connection>
<GID>589</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,-11,196.5,-11</points>
<connection>
<GID>590</GID>
<name>IN_0</name></connection>
<intersection>195 0</intersection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213.5,-11,213.5,-9</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213.5,-11,215,-11</points>
<connection>
<GID>598</GID>
<name>IN_0</name></connection>
<intersection>213.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-11,222.5,-9</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-11,224,-11</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-11,231.5,-9</points>
<connection>
<GID>605</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,-11,233,-11</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<intersection>231.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>574</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240.5,-11,240.5,-9</points>
<connection>
<GID>609</GID>
<name>OUT</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240.5,-11,242,-11</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>240.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,3,241.5,13.5</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,13.5,241.5,13.5</points>
<connection>
<GID>613</GID>
<name>OUT_7</name></connection>
<intersection>241.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,3,232.5,12.5</points>
<connection>
<GID>604</GID>
<name>IN_1</name></connection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,12.5,232.5,12.5</points>
<connection>
<GID>613</GID>
<name>OUT_6</name></connection>
<intersection>232.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223.5,3,223.5,11.5</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,11.5,223.5,11.5</points>
<connection>
<GID>613</GID>
<name>OUT_5</name></connection>
<intersection>223.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,3,214.5,10.5</points>
<connection>
<GID>596</GID>
<name>IN_1</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,10.5,214.5,10.5</points>
<connection>
<GID>613</GID>
<name>OUT_4</name></connection>
<intersection>214.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,3,205,9.5</points>
<connection>
<GID>592</GID>
<name>IN_1</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,9.5,205,9.5</points>
<connection>
<GID>613</GID>
<name>OUT_3</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>580</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,3,196,8.5</points>
<connection>
<GID>588</GID>
<name>IN_1</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,8.5,196,8.5</points>
<connection>
<GID>613</GID>
<name>OUT_2</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>581</ID>
<shape>
<hsegment>
<ID>58</ID>
<points>181,-44.5,436,-44.5</points>
<connection>
<GID>656</GID>
<name>OUT</name></connection>
<intersection>366.5 148</intersection>
<intersection>372.5 1066</intersection>
<intersection>381.5 1067</intersection>
<intersection>390.5 1065</intersection>
<intersection>400 1068</intersection>
<intersection>409 1064</intersection>
<intersection>418 1069</intersection>
<intersection>427 1063</intersection>
<intersection>436 1070</intersection></hsegment>
<vsegment>
<ID>148</ID>
<points>366.5,-97,366.5,-44.5</points>
<intersection>-97 150</intersection>
<intersection>-44.5 58</intersection></vsegment>
<hsegment>
<ID>150</ID>
<points>366.5,-97,437.5,-97</points>
<intersection>366.5 148</intersection>
<intersection>374 1019</intersection>
<intersection>383 1060</intersection>
<intersection>392 1058</intersection>
<intersection>401.5 1061</intersection>
<intersection>410.5 1057</intersection>
<intersection>419.5 1062</intersection>
<intersection>428.5 1056</intersection>
<intersection>437.5 180</intersection></hsegment>
<vsegment>
<ID>180</ID>
<points>437.5,-123,437.5,-86</points>
<connection>
<GID>695</GID>
<name>clock</name></connection>
<intersection>-123 1042</intersection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1019</ID>
<points>374,-97,374,-86</points>
<connection>
<GID>665</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<hsegment>
<ID>1042</ID>
<points>437.5,-123,560,-123</points>
<intersection>437.5 180</intersection>
<intersection>560 1043</intersection></hsegment>
<vsegment>
<ID>1043</ID>
<points>560,-123,560,-109</points>
<intersection>-123 1042</intersection>
<intersection>-109 1046</intersection></vsegment>
<hsegment>
<ID>1046</ID>
<points>560,-109,564.5,-109</points>
<connection>
<GID>810</GID>
<name>IN_1</name></connection>
<intersection>560 1043</intersection></hsegment>
<vsegment>
<ID>1056</ID>
<points>428.5,-97,428.5,-86</points>
<connection>
<GID>691</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1057</ID>
<points>410.5,-97,410.5,-86</points>
<connection>
<GID>683</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1058</ID>
<points>392,-97,392,-86</points>
<connection>
<GID>675</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1060</ID>
<points>383,-97,383,-86</points>
<connection>
<GID>671</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1061</ID>
<points>401.5,-97,401.5,-86</points>
<connection>
<GID>679</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1062</ID>
<points>419.5,-97,419.5,-86</points>
<connection>
<GID>687</GID>
<name>clock</name></connection>
<intersection>-97 150</intersection></vsegment>
<vsegment>
<ID>1063</ID>
<points>427,-44.5,427,-26.5</points>
<connection>
<GID>727</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1064</ID>
<points>409,-44.5,409,-26.5</points>
<connection>
<GID>719</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1065</ID>
<points>390.5,-44.5,390.5,-26.5</points>
<connection>
<GID>711</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1066</ID>
<points>372.5,-44.5,372.5,-26.5</points>
<connection>
<GID>700</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1067</ID>
<points>381.5,-44.5,381.5,-26.5</points>
<connection>
<GID>706</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1068</ID>
<points>400,-44.5,400,-26.5</points>
<connection>
<GID>715</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1069</ID>
<points>418,-44.5,418,-26.5</points>
<connection>
<GID>723</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment>
<vsegment>
<ID>1070</ID>
<points>436,-44.5,436,-26.5</points>
<connection>
<GID>731</GID>
<name>clock</name></connection>
<intersection>-44.5 58</intersection></vsegment></shape></wire>
<wire>
<ID>582</ID>
<shape>
<vsegment>
<ID>11</ID>
<points>155,-37,155,-35.5</points>
<connection>
<GID>616</GID>
<name>IN_1</name></connection>
<connection>
<GID>615</GID>
<name>CLK</name></connection></vsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-31.5,148.5,-31.5</points>
<connection>
<GID>619</GID>
<name>OUT_0</name></connection>
<connection>
<GID>620</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>584</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-33.5,155,-32.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>-32.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>154.5,-32.5,155,-32.5</points>
<connection>
<GID>620</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141,-33.5,148.5,-33.5</points>
<connection>
<GID>620</GID>
<name>IN_1</name></connection>
<intersection>141 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>141,-40,141,-28</points>
<connection>
<GID>582</GID>
<name>OUT_0</name></connection>
<intersection>-40 16</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>141,-40,153.5,-40</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>141 9</intersection></hsegment></shape></wire>
<wire>
<ID>586</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>164.5,-40,164.5,-33.5</points>
<connection>
<GID>583</GID>
<name>IN_1</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-40,164.5,-40</points>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection>
<intersection>164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160.5,-27.5,163.5,-27.5</points>
<connection>
<GID>583</GID>
<name>OUT</name></connection>
<connection>
<GID>617</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-26.5,151.5,-26.5</points>
<connection>
<GID>617</GID>
<name>count_enable</name></connection>
<connection>
<GID>618</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-31.5,144.5,-15.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-15.5,163.5,-15.5</points>
<intersection>144.5 0</intersection>
<intersection>156 3</intersection>
<intersection>163.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>163.5,-25.5,163.5,-15.5</points>
<intersection>-25.5 4</intersection>
<intersection>-15.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>156,-16,156,-15.5</points>
<connection>
<GID>550</GID>
<name>OUT</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>160.5,-25.5,163.5,-25.5</points>
<connection>
<GID>617</GID>
<name>clear</name></connection>
<intersection>163.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-22.5,154.5,-22</points>
<connection>
<GID>617</GID>
<name>OUT_3</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>154.5,-22,155,-22</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-25.5,309,-21</points>
<connection>
<GID>622</GID>
<name>OUT_0</name></connection>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,-21,332,-21</points>
<intersection>309 0</intersection>
<intersection>332 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>332,-21,332,-5.5</points>
<intersection>-21 1</intersection>
<intersection>-5.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>332,-5.5,334,-5.5</points>
<connection>
<GID>621</GID>
<name>IN_0</name></connection>
<intersection>332 2</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-17,309,-12</points>
<connection>
<GID>623</GID>
<name>OUT_0</name></connection>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,-12,331,-12</points>
<intersection>309 0</intersection>
<intersection>331 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>331,-12,331,-4.5</points>
<intersection>-12 3</intersection>
<intersection>-4.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>331,-4.5,334,-4.5</points>
<connection>
<GID>621</GID>
<name>IN_1</name></connection>
<intersection>331 4</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-8.5,309,-3.5</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<intersection>-3.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>309,-3.5,334,-3.5</points>
<connection>
<GID>621</GID>
<name>IN_2</name></connection>
<intersection>309 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-0.5,309,4.5</points>
<connection>
<GID>625</GID>
<name>OUT_0</name></connection>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,4.5,329,4.5</points>
<intersection>309 0</intersection>
<intersection>329 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>329,-2.5,329,4.5</points>
<intersection>-2.5 5</intersection>
<intersection>4.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>329,-2.5,334,-2.5</points>
<connection>
<GID>621</GID>
<name>IN_3</name></connection>
<intersection>329 4</intersection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>330,-1.5,330,8</points>
<intersection>-1.5 5</intersection>
<intersection>8 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>330,-1.5,334,-1.5</points>
<connection>
<GID>621</GID>
<name>IN_4</name></connection>
<intersection>330 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>309,8,330,8</points>
<intersection>309 8</intersection>
<intersection>330 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>309,7,309,8.5</points>
<connection>
<GID>626</GID>
<name>OUT_0</name></connection>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>8 6</intersection></vsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,14.5,309,19.5</points>
<connection>
<GID>627</GID>
<name>OUT_0</name></connection>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>19.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,19.5,331,19.5</points>
<intersection>309 0</intersection>
<intersection>331 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>331,-0.5,331,19.5</points>
<intersection>-0.5 5</intersection>
<intersection>19.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>331,-0.5,334,-0.5</points>
<connection>
<GID>621</GID>
<name>IN_5</name></connection>
<intersection>331 4</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,22,309,27</points>
<connection>
<GID>628</GID>
<name>OUT_0</name></connection>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>309,27,332,27</points>
<intersection>309 0</intersection>
<intersection>332 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>332,0.5,332,27</points>
<intersection>0.5 5</intersection>
<intersection>27 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>332,0.5,334,0.5</points>
<connection>
<GID>621</GID>
<name>IN_6</name></connection>
<intersection>332 4</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,29.5,309,30</points>
<connection>
<GID>629</GID>
<name>OUT_0</name></connection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309,30,334,30</points>
<intersection>309 0</intersection>
<intersection>334 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>334,1.5,334,30</points>
<connection>
<GID>621</GID>
<name>IN_7</name></connection>
<intersection>30 1</intersection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>337,3.5,337,3.5</points>
<connection>
<GID>621</GID>
<name>load</name></connection>
<connection>
<GID>631</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-108.5,311,-106</points>
<connection>
<GID>633</GID>
<name>OUT_0</name></connection>
<connection>
<GID>634</GID>
<name>IN_0</name></connection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-107,334,-107</points>
<intersection>311 0</intersection>
<intersection>334 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>334,-107,334,-88.5</points>
<intersection>-107 1</intersection>
<intersection>-88.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>334,-88.5,336,-88.5</points>
<connection>
<GID>632</GID>
<name>IN_0</name></connection>
<intersection>334 2</intersection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-100,311,-98</points>
<connection>
<GID>634</GID>
<name>OUT_0</name></connection>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<intersection>-99 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>311,-99,333,-99</points>
<intersection>311 0</intersection>
<intersection>333 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>333,-99,333,-87.5</points>
<intersection>-99 3</intersection>
<intersection>-87.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>333,-87.5,336,-87.5</points>
<connection>
<GID>632</GID>
<name>IN_1</name></connection>
<intersection>333 4</intersection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-92,311,-90</points>
<connection>
<GID>635</GID>
<name>OUT_0</name></connection>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<intersection>-91 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>311,-91,336,-91</points>
<intersection>311 0</intersection>
<intersection>336 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>336,-91,336,-86.5</points>
<connection>
<GID>632</GID>
<name>IN_2</name></connection>
<intersection>-91 6</intersection></vsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-84,311,-82</points>
<connection>
<GID>636</GID>
<name>OUT_0</name></connection>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>311,-83,331,-83</points>
<intersection>311 0</intersection>
<intersection>331 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>331,-85.5,331,-83</points>
<intersection>-85.5 5</intersection>
<intersection>-83 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>331,-85.5,336,-85.5</points>
<connection>
<GID>632</GID>
<name>IN_3</name></connection>
<intersection>331 4</intersection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,-84.5,332,-75</points>
<intersection>-84.5 5</intersection>
<intersection>-75 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>332,-84.5,336,-84.5</points>
<connection>
<GID>632</GID>
<name>IN_4</name></connection>
<intersection>332 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>311,-75,332,-75</points>
<intersection>311 8</intersection>
<intersection>332 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>311,-76,311,-74</points>
<connection>
<GID>637</GID>
<name>OUT_0</name></connection>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>-75 6</intersection></vsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-68,311,-66</points>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection>
<connection>
<GID>639</GID>
<name>IN_0</name></connection>
<intersection>-67 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>311,-67,333,-67</points>
<intersection>311 0</intersection>
<intersection>333 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>333,-83.5,333,-67</points>
<intersection>-83.5 5</intersection>
<intersection>-67 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>333,-83.5,336,-83.5</points>
<connection>
<GID>632</GID>
<name>IN_5</name></connection>
<intersection>333 4</intersection></hsegment></shape></wire>
<wire>
<ID>609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-60,311,-58</points>
<connection>
<GID>639</GID>
<name>OUT_0</name></connection>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>311,-59,334,-59</points>
<intersection>311 0</intersection>
<intersection>334 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>334,-82.5,334,-59</points>
<intersection>-82.5 5</intersection>
<intersection>-59 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>334,-82.5,336,-82.5</points>
<connection>
<GID>632</GID>
<name>IN_6</name></connection>
<intersection>334 4</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311,-52,311,-51</points>
<connection>
<GID>640</GID>
<name>OUT_0</name></connection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311,-51,336,-51</points>
<intersection>311 0</intersection>
<intersection>336 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>336,-81.5,336,-51</points>
<connection>
<GID>632</GID>
<name>IN_7</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156.5,-14.5,172,-14.5</points>
<intersection>156.5 7</intersection>
<intersection>172 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>172,-31.5,172,-14.5</points>
<intersection>-31.5 5</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>172,-31.5,184.5,-31.5</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<intersection>172 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>156.5,-14.5,156.5,-12</points>
<intersection>-14.5 1</intersection>
<intersection>-12 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>154.5,-12,157.5,-12</points>
<connection>
<GID>815</GID>
<name>OUT</name></connection>
<connection>
<GID>641</GID>
<name>IN_1</name></connection>
<intersection>156.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>339,-79.5,339,-79.5</points>
<connection>
<GID>632</GID>
<name>load</name></connection>
<connection>
<GID>642</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,13.5,158.5,15.5</points>
<intersection>13.5 1</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,13.5,164.5,13.5</points>
<connection>
<GID>613</GID>
<name>IN_7</name></connection>
<intersection>158.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,15.5,158.5,15.5</points>
<connection>
<GID>643</GID>
<name>OUT_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,12.5,157.5,13.5</points>
<intersection>12.5 2</intersection>
<intersection>13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,13.5,157.5,13.5</points>
<connection>
<GID>644</GID>
<name>OUT_0</name></connection>
<intersection>157.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,12.5,164.5,12.5</points>
<connection>
<GID>613</GID>
<name>IN_6</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>143.5,11.5,164.5,11.5</points>
<connection>
<GID>613</GID>
<name>IN_5</name></connection>
<connection>
<GID>645</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,9.5,157,10.5</points>
<intersection>9.5 1</intersection>
<intersection>10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,9.5,157,9.5</points>
<connection>
<GID>646</GID>
<name>OUT_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,10.5,164.5,10.5</points>
<connection>
<GID>613</GID>
<name>IN_4</name></connection>
<intersection>157 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,7.5,158,9.5</points>
<intersection>7.5 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,9.5,164.5,9.5</points>
<connection>
<GID>613</GID>
<name>IN_3</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,7.5,158,7.5</points>
<connection>
<GID>647</GID>
<name>OUT_0</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>143.5,5.5,159,5.5</points>
<connection>
<GID>648</GID>
<name>OUT_0</name></connection>
<intersection>159 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>159,5.5,159,8.5</points>
<intersection>5.5 1</intersection>
<intersection>8.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>159,8.5,164.5,8.5</points>
<connection>
<GID>613</GID>
<name>IN_2</name></connection>
<intersection>159 3</intersection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,1.5,161,6.5</points>
<intersection>1.5 2</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,6.5,164.5,6.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,1.5,161,1.5</points>
<connection>
<GID>650</GID>
<name>OUT_0</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,3.5,160,7.5</points>
<intersection>3.5 1</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,3.5,160,3.5</points>
<connection>
<GID>649</GID>
<name>OUT_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,7.5,164.5,7.5</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,15.5,167.5,15.5</points>
<connection>
<GID>613</GID>
<name>load</name></connection>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-22.5,157.5,-22</points>
<connection>
<GID>617</GID>
<name>OUT_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>157,-22,157.5,-22</points>
<connection>
<GID>550</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-11,163.5,-3.5</points>
<connection>
<GID>641</GID>
<name>OUT</name></connection>
<connection>
<GID>816</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>456.5,-70.5,560.5,-70.5</points>
<connection>
<GID>661</GID>
<name>IN_1</name></connection>
<intersection>456.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>456.5,-70.5,456.5,-57.5</points>
<connection>
<GID>660</GID>
<name>OUT</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>626</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>174.5,-43.5,174.5,-37</points>
<intersection>-43.5 6</intersection>
<intersection>-37 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>173,-37,175,-37</points>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<intersection>174.5 1</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>174.5,-43.5,175,-43.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<intersection>174.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>379.5,-75,380.5,-75</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<connection>
<GID>666</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>628</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>382.5,-75,383.5,-75</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<connection>
<GID>667</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>629</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-10,154,25</points>
<intersection>-10 10</intersection>
<intersection>-7.5 5</intersection>
<intersection>-3.5 13</intersection>
<intersection>25 19</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>154,-7.5,175,-7.5</points>
<intersection>154 0</intersection>
<intersection>175 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>175,-35,175,-7.5</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-7.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>154,-10,157.5,-10</points>
<connection>
<GID>641</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>152,-3.5,154,-3.5</points>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>153.5,25,154,25</points>
<connection>
<GID>813</GID>
<name>OUT_0</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>630</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>377,-80.5,377,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>377,-80.5,380,-80.5</points>
<intersection>377 0</intersection>
<intersection>380 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>377,-69,378.5,-69</points>
<connection>
<GID>666</GID>
<name>IN_1</name></connection>
<intersection>377 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>380,-83,380,-80.5</points>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>631</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>388.5,-75,389.5,-75</points>
<connection>
<GID>674</GID>
<name>IN_1</name></connection>
<connection>
<GID>672</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>632</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>391.5,-75,392.5,-75</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<connection>
<GID>673</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>633</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386,-80.5,386,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>386,-80.5,389,-80.5</points>
<intersection>386 0</intersection>
<intersection>389 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>386,-69,387.5,-69</points>
<connection>
<GID>672</GID>
<name>IN_1</name></connection>
<intersection>386 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>389,-83,389,-80.5</points>
<connection>
<GID>671</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>634</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>397.5,-75,398.5,-75</points>
<connection>
<GID>678</GID>
<name>IN_1</name></connection>
<connection>
<GID>676</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>635</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>400.5,-75,401.5,-75</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<connection>
<GID>677</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>395,-80.5,395,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>395,-80.5,398,-80.5</points>
<intersection>395 0</intersection>
<intersection>398 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>395,-69,396.5,-69</points>
<connection>
<GID>676</GID>
<name>IN_1</name></connection>
<intersection>395 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>398,-83,398,-80.5</points>
<connection>
<GID>675</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>407,-75,408,-75</points>
<connection>
<GID>682</GID>
<name>IN_1</name></connection>
<connection>
<GID>680</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>638</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>410,-75,411,-75</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<connection>
<GID>681</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>404.5,-80.5,404.5,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>404.5,-80.5,407.5,-80.5</points>
<intersection>404.5 0</intersection>
<intersection>407.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>404.5,-69,406,-69</points>
<connection>
<GID>680</GID>
<name>IN_1</name></connection>
<intersection>404.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>407.5,-83,407.5,-80.5</points>
<connection>
<GID>679</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>416,-75,417,-75</points>
<connection>
<GID>686</GID>
<name>IN_1</name></connection>
<connection>
<GID>684</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>641</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>419,-75,420,-75</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<connection>
<GID>685</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>413.5,-80.5,413.5,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>413.5,-80.5,416.5,-80.5</points>
<intersection>413.5 0</intersection>
<intersection>416.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>413.5,-69,415,-69</points>
<connection>
<GID>684</GID>
<name>IN_1</name></connection>
<intersection>413.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>416.5,-83,416.5,-80.5</points>
<connection>
<GID>683</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>425,-75,426,-75</points>
<connection>
<GID>690</GID>
<name>IN_1</name></connection>
<connection>
<GID>688</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>644</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>428,-75,429,-75</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<connection>
<GID>689</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,-80.5,422.5,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>422.5,-80.5,425.5,-80.5</points>
<intersection>422.5 0</intersection>
<intersection>425.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,-69,424,-69</points>
<connection>
<GID>688</GID>
<name>IN_1</name></connection>
<intersection>422.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>425.5,-83,425.5,-80.5</points>
<connection>
<GID>687</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>646</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>434,-75,435,-75</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<connection>
<GID>692</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>437,-75,438,-75</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>431.5,-80.5,431.5,-69</points>
<intersection>-80.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>431.5,-80.5,434.5,-80.5</points>
<intersection>431.5 0</intersection>
<intersection>434.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>431.5,-69,433,-69</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<intersection>431.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>434.5,-83,434.5,-80.5</points>
<connection>
<GID>691</GID>
<name>OUT_0</name></connection>
<intersection>-80.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>161,-34.5,166,-34.5</points>
<connection>
<GID>616</GID>
<name>OUT</name></connection>
<intersection>162.5 10</intersection>
<intersection>166 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>166,-38,166,-34.5</points>
<intersection>-38 9</intersection>
<intersection>-36 8</intersection>
<intersection>-34.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>166,-36,167,-36</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<intersection>166 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>166,-38,167,-38</points>
<connection>
<GID>571</GID>
<name>IN_1</name></connection>
<intersection>166 7</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>162.5,-34.5,162.5,-33.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<intersection>-34.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-18.5,178.5,-14</points>
<connection>
<GID>577</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-18.5,242,-18.5</points>
<intersection>178.5 0</intersection>
<intersection>181 3</intersection>
<intersection>187.5 10</intersection>
<intersection>196.5 9</intersection>
<intersection>206 8</intersection>
<intersection>215 7</intersection>
<intersection>224 6</intersection>
<intersection>233 5</intersection>
<intersection>242 41</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>181,-36,181,-18.5</points>
<connection>
<GID>653</GID>
<name>OUT</name></connection>
<intersection>-36 12</intersection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>233,-18.5,233,-14</points>
<connection>
<GID>606</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>224,-18.5,224,-14</points>
<connection>
<GID>602</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>215,-18.5,215,-14</points>
<connection>
<GID>598</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>206,-18.5,206,-14</points>
<connection>
<GID>594</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>196.5,-18.5,196.5,-14</points>
<connection>
<GID>590</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>187.5,-18.5,187.5,-14</points>
<connection>
<GID>585</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>181,-36,258.5,-36</points>
<intersection>181 3</intersection>
<intersection>258.5 36</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>258.5,-55.5,258.5,-36</points>
<intersection>-55.5 38</intersection>
<intersection>-47.5 39</intersection>
<intersection>-36 12</intersection></vsegment>
<hsegment>
<ID>38</ID>
<points>258.5,-55.5,278.5,-55.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>258.5 36</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>258.5,-47.5,278.5,-47.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<intersection>258.5 36</intersection></hsegment>
<vsegment>
<ID>41</ID>
<points>242,-18.5,242,-14</points>
<connection>
<GID>611</GID>
<name>clock</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>381.5,-83,381.5,-81</points>
<connection>
<GID>668</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>381.5,-83,383,-83</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>381.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399.5,-83,399.5,-81</points>
<connection>
<GID>678</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>399.5,-83,401.5,-83</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>399.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>390.5,-83,390.5,-81</points>
<connection>
<GID>674</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>390.5,-83,392,-83</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>390.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>409,-83,409,-81</points>
<connection>
<GID>682</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>409,-83,410.5,-83</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>409 0</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418,-83,418,-81</points>
<connection>
<GID>686</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418,-83,419.5,-83</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>418 0</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427,-83,427,-81</points>
<connection>
<GID>690</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427,-83,428.5,-83</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>427 0</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,-83,436,-81</points>
<connection>
<GID>694</GID>
<name>OUT</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436,-83,437.5,-83</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>436 0</intersection></hsegment></shape></wire>
<wire>
<ID>658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-31.5,201,-27</points>
<intersection>-31.5 16</intersection>
<intersection>-30.5 8</intersection>
<intersection>-29.5 7</intersection>
<intersection>-27 18</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>201,-29.5,202,-29.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>200.5,-30.5,201,-30.5</points>
<connection>
<GID>670</GID>
<name>OUT_0</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>201,-31.5,202,-31.5</points>
<connection>
<GID>669</GID>
<name>IN_1</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>201,-27,202,-27</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>141,-24,141,-24</points>
<connection>
<GID>579</GID>
<name>OUT_0</name></connection>
<connection>
<GID>582</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180.5,3.5,243.5,3.5</points>
<connection>
<GID>584</GID>
<name>OUT_0</name></connection>
<intersection>189 4</intersection>
<intersection>198 6</intersection>
<intersection>207 7</intersection>
<intersection>216.5 8</intersection>
<intersection>225.5 9</intersection>
<intersection>234.5 10</intersection>
<intersection>243.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243.5,3,243.5,3.5</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>189,3,189,3.5</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>198,3,198,3.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>207,3,207,3.5</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>216.5,3,216.5,3.5</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>225.5,3,225.5,3.5</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>234.5,3,234.5,3.5</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190.5,-30.5,196.5,-30.5</points>
<connection>
<GID>657</GID>
<name>OUT</name></connection>
<connection>
<GID>670</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,3,185,5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174.5,5,239.5,5</points>
<intersection>174.5 2</intersection>
<intersection>185 0</intersection>
<intersection>194 5</intersection>
<intersection>203 6</intersection>
<intersection>212.5 7</intersection>
<intersection>221.5 8</intersection>
<intersection>230.5 9</intersection>
<intersection>239.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>174.5,-2.5,174.5,5</points>
<connection>
<GID>698</GID>
<name>OUT</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>239.5,3,239.5,5</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>194,3,194,5</points>
<connection>
<GID>587</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>203,3,203,5</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>212.5,3,212.5,5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>221.5,3,221.5,5</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>230.5,3,230.5,5</points>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment></shape></wire>
<wire>
<ID>665</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>164.5,4.5,167.5,4.5</points>
<connection>
<GID>696</GID>
<name>CLK</name></connection>
<connection>
<GID>613</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>378,-15.5,379,-15.5</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<connection>
<GID>701</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>667</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>381,-15.5,382,-15.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<connection>
<GID>703</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>668</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>456,-116.5,458.5,-116.5</points>
<connection>
<GID>736</GID>
<name>IN_1</name></connection>
<intersection>456 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>456,-117.5,456,-116.5</points>
<intersection>-117.5 12</intersection>
<intersection>-116.5 3</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>453,-117.5,456,-117.5</points>
<connection>
<GID>735</GID>
<name>CLK</name></connection>
<intersection>456 11</intersection></hsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-112.5,452,-112.5</points>
<connection>
<GID>739</GID>
<name>OUT_0</name></connection>
<connection>
<GID>740</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375.5,-21,375.5,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375.5,-21,378.5,-21</points>
<intersection>375.5 0</intersection>
<intersection>378.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>375.5,-9.5,377,-9.5</points>
<connection>
<GID>701</GID>
<name>IN_1</name></connection>
<intersection>375.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>378.5,-23.5,378.5,-21</points>
<connection>
<GID>700</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>671</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>387,-15.5,388,-15.5</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<connection>
<GID>708</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>672</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>390,-15.5,391,-15.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<connection>
<GID>709</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-21,384.5,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-21,387.5,-21</points>
<intersection>384.5 0</intersection>
<intersection>387.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>384.5,-9.5,386,-9.5</points>
<connection>
<GID>708</GID>
<name>IN_1</name></connection>
<intersection>384.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>387.5,-23.5,387.5,-21</points>
<connection>
<GID>706</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>674</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>396,-15.5,397,-15.5</points>
<connection>
<GID>714</GID>
<name>IN_1</name></connection>
<connection>
<GID>712</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>675</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>399,-15.5,400,-15.5</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<connection>
<GID>713</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393.5,-21,393.5,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>393.5,-21,396.5,-21</points>
<intersection>393.5 0</intersection>
<intersection>396.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>393.5,-9.5,395,-9.5</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>393.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>396.5,-23.5,396.5,-21</points>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>677</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>405.5,-15.5,406.5,-15.5</points>
<connection>
<GID>718</GID>
<name>IN_1</name></connection>
<connection>
<GID>716</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>678</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>408.5,-15.5,409.5,-15.5</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<connection>
<GID>717</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>403,-21,403,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403,-21,406,-21</points>
<intersection>403 0</intersection>
<intersection>406 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403,-9.5,404.5,-9.5</points>
<connection>
<GID>716</GID>
<name>IN_1</name></connection>
<intersection>403 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>406,-23.5,406,-21</points>
<connection>
<GID>715</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>680</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>414.5,-15.5,415.5,-15.5</points>
<connection>
<GID>722</GID>
<name>IN_1</name></connection>
<connection>
<GID>720</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>681</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>417.5,-15.5,418.5,-15.5</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<connection>
<GID>721</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,-21,412,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>412,-21,415,-21</points>
<intersection>412 0</intersection>
<intersection>415 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,-9.5,413.5,-9.5</points>
<connection>
<GID>720</GID>
<name>IN_1</name></connection>
<intersection>412 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>415,-23.5,415,-21</points>
<connection>
<GID>719</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>683</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>423.5,-15.5,424.5,-15.5</points>
<connection>
<GID>726</GID>
<name>IN_1</name></connection>
<connection>
<GID>724</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>684</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>426.5,-15.5,427.5,-15.5</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<connection>
<GID>725</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421,-21,421,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>421,-21,424,-21</points>
<intersection>421 0</intersection>
<intersection>424 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421,-9.5,422.5,-9.5</points>
<connection>
<GID>724</GID>
<name>IN_1</name></connection>
<intersection>421 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>424,-23.5,424,-21</points>
<connection>
<GID>723</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>432.5,-15.5,433.5,-15.5</points>
<connection>
<GID>730</GID>
<name>IN_1</name></connection>
<connection>
<GID>728</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>687</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>435.5,-15.5,436.5,-15.5</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<connection>
<GID>729</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>430,-21,430,-9.5</points>
<intersection>-21 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>430,-21,433,-21</points>
<intersection>430 0</intersection>
<intersection>433 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>430,-9.5,431.5,-9.5</points>
<connection>
<GID>728</GID>
<name>IN_1</name></connection>
<intersection>430 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>433,-23.5,433,-21</points>
<connection>
<GID>727</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>458.5,-114.5,458.5,-113.5</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<intersection>-113.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>458,-113.5,458.5,-113.5</points>
<connection>
<GID>740</GID>
<name>OUT</name></connection>
<intersection>458.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>444.5,-114.5,452,-114.5</points>
<connection>
<GID>740</GID>
<name>IN_1</name></connection>
<intersection>444.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>444.5,-120,444.5,-109</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>-120 16</intersection>
<intersection>-114.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>444.5,-120,457,-120</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<intersection>444.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-23.5,380,-21.5</points>
<connection>
<GID>704</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-23.5,381.5,-23.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-23.5,398,-21.5</points>
<connection>
<GID>714</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,-23.5,400,-23.5</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<intersection>398 0</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-23.5,389,-21.5</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>389,-23.5,390.5,-23.5</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>389 0</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>407.5,-23.5,407.5,-21.5</points>
<connection>
<GID>718</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>407.5,-23.5,409,-23.5</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>407.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416.5,-23.5,416.5,-21.5</points>
<connection>
<GID>722</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>416.5,-23.5,418,-23.5</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<intersection>416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>425.5,-23.5,425.5,-21.5</points>
<connection>
<GID>726</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>425.5,-23.5,427,-23.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<intersection>425.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-23.5,434.5,-21.5</points>
<connection>
<GID>730</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,-23.5,436,-23.5</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,-120,468,-114.5</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>461,-120,468,-120</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>468 0</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>464,-108.5,467,-108.5</points>
<connection>
<GID>733</GID>
<name>OUT</name></connection>
<connection>
<GID>737</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-3.5,168.5,3.5</points>
<connection>
<GID>698</GID>
<name>IN_1</name></connection>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>-3.5 8</intersection>
<intersection>3.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>168.5,3.5,176.5,3.5</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>167.5,-3.5,168.5,-3.5</points>
<connection>
<GID>816</GID>
<name>OUT_0</name></connection>
<intersection>168.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455,-107.5,455,-107.5</points>
<connection>
<GID>737</GID>
<name>count_enable</name></connection>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,-112.5,448,-97</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>448,-97,467,-97</points>
<connection>
<GID>702</GID>
<name>OUT</name></connection>
<intersection>448 0</intersection>
<intersection>467 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>467,-106.5,467,-97</points>
<intersection>-106.5 4</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>464,-106.5,467,-106.5</points>
<connection>
<GID>737</GID>
<name>clear</name></connection>
<intersection>467 2</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>458,-103,458.5,-103</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>458 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>458,-103.5,458,-103</points>
<connection>
<GID>737</GID>
<name>OUT_3</name></connection>
<intersection>-103 2</intersection></vsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>460.5,-103,461,-103</points>
<connection>
<GID>702</GID>
<name>IN_1</name></connection>
<intersection>461 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>461,-103.5,461,-103</points>
<connection>
<GID>737</GID>
<name>OUT_0</name></connection>
<intersection>-103 2</intersection></vsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>463.5,-92.5,466,-92.5</points>
<connection>
<GID>797</GID>
<name>IN_0</name></connection>
<intersection>463.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>463.5,-93.5,463.5,-92.5</points>
<intersection>-93.5 11</intersection>
<intersection>-92.5 5</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>458,-93.5,463.5,-93.5</points>
<connection>
<GID>796</GID>
<name>OUT</name></connection>
<intersection>463.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>464.5,-115.5,471.5,-115.5</points>
<connection>
<GID>736</GID>
<name>OUT</name></connection>
<intersection>466 34</intersection>
<intersection>471.5 37</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>466,-115.5,466,-114.5</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>-115.5 6</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>471.5,-116.5,471.5,-114.5</points>
<connection>
<GID>705</GID>
<name>IN_1</name></connection>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>-115.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>444.5,-105,444.5,-105</points>
<connection>
<GID>707</GID>
<name>OUT_0</name></connection>
<connection>
<GID>732</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-96.5,470,-92.5</points>
<connection>
<GID>797</GID>
<name>OUT_0</name></connection>
<intersection>-96.5 27</intersection>
<intersection>-92.5 29</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>470,-96.5,478.5,-96.5</points>
<intersection>470 0</intersection>
<intersection>478.5 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>478.5,-96.5,478.5,-85.5</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>-96.5 27</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>470,-92.5,471,-92.5</points>
<intersection>470 0</intersection>
<intersection>471 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>471,-93.5,471,-91.5</points>
<connection>
<GID>747</GID>
<name>IN_1</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>-92.5 29</intersection></vsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>444.5,-101,444.5,-94.5</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>-94.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>444.5,-94.5,448,-94.5</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<intersection>444.5 7</intersection>
<intersection>448 28</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>448,-94.5,448,-82.5</points>
<intersection>-94.5 10</intersection>
<intersection>-92.5 29</intersection>
<intersection>-82.5 45</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>448,-92.5,452,-92.5</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<intersection>448 28</intersection></hsegment>
<hsegment>
<ID>45</ID>
<points>448,-82.5,453,-82.5</points>
<connection>
<GID>809</GID>
<name>OUT_0</name></connection>
<intersection>448 28</intersection></hsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452,-94.5,452,-94.5</points>
<connection>
<GID>773</GID>
<name>OUT_0</name></connection>
<connection>
<GID>796</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-101.5,277.5,33</points>
<connection>
<GID>576</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 13</intersection>
<intersection>-85.5 10</intersection>
<intersection>-69.5 5</intersection>
<intersection>-53.5 1</intersection>
<intersection>-27 28</intersection>
<intersection>-11 25</intersection>
<intersection>5 20</intersection>
<intersection>21 16</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277.5,-53.5,278.5,-53.5</points>
<connection>
<GID>575</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>277.5,-69.5,278.5,-69.5</points>
<connection>
<GID>630</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>277.5,-85.5,278.5,-85.5</points>
<connection>
<GID>699</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>277.5,-101.5,278.5,-101.5</points>
<connection>
<GID>800</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>277.5,21,278.5,21</points>
<connection>
<GID>556</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>277.5,5,278.5,5</points>
<connection>
<GID>560</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>277.5,-11,278.5,-11</points>
<connection>
<GID>564</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>277.5,-27,278.5,-27</points>
<connection>
<GID>568</GID>
<name>IN_3</name></connection>
<intersection>277.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>477.5,-107.5,557.5,-107.5</points>
<intersection>477.5 20</intersection>
<intersection>481.5 9</intersection>
<intersection>491.5 8</intersection>
<intersection>501.5 7</intersection>
<intersection>511.5 6</intersection>
<intersection>521.5 16</intersection>
<intersection>531.5 12</intersection>
<intersection>541.5 14</intersection>
<intersection>551.5 11</intersection>
<intersection>557.5 24</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>511.5,-107.5,511.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>501.5,-107.5,501.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>491.5,-107.5,491.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>481.5,-107.5,481.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>551.5,-107.5,551.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>531.5,-107.5,531.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>541.5,-107.5,541.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>521.5,-107.5,521.5,-103.5</points>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>477.5,-115.5,477.5,-103.5</points>
<connection>
<GID>705</GID>
<name>OUT</name></connection>
<intersection>-107.5 2</intersection>
<intersection>-103.5 28</intersection></vsegment>
<vsegment>
<ID>24</ID>
<points>557.5,-107.5,557.5,-107</points>
<intersection>-107.5 2</intersection>
<intersection>-107 25</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>557.5,-107,564.5,-107</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<intersection>557.5 24</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>477.5,-103.5,552.5,-103.5</points>
<connection>
<GID>772</GID>
<name>clock</name></connection>
<connection>
<GID>742</GID>
<name>clock</name></connection>
<connection>
<GID>748</GID>
<name>clock</name></connection>
<connection>
<GID>752</GID>
<name>clock</name></connection>
<connection>
<GID>756</GID>
<name>clock</name></connection>
<connection>
<GID>760</GID>
<name>clock</name></connection>
<connection>
<GID>764</GID>
<name>clock</name></connection>
<connection>
<GID>768</GID>
<name>clock</name></connection>
<intersection>477.5 20</intersection>
<intersection>481.5 9</intersection>
<intersection>491.5 8</intersection>
<intersection>501.5 7</intersection>
<intersection>511.5 6</intersection>
<intersection>521.5 16</intersection>
<intersection>531.5 12</intersection>
<intersection>541.5 14</intersection>
<intersection>551.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>488.5,-92.5,489.5,-92.5</points>
<connection>
<GID>745</GID>
<name>IN_1</name></connection>
<connection>
<GID>743</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>491.5,-92.5,492.5,-92.5</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<connection>
<GID>744</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-84,549.5,-84</points>
<intersection>477.5 27</intersection>
<intersection>489.5 42</intersection>
<intersection>499.5 34</intersection>
<intersection>509.5 37</intersection>
<intersection>519.5 38</intersection>
<intersection>529.5 39</intersection>
<intersection>539.5 40</intersection>
<intersection>549.5 36</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>477.5,-92.5,477.5,-84</points>
<intersection>-92.5 43</intersection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>34</ID>
<points>499.5,-86.5,499.5,-84</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>549.5,-86.5,549.5,-84</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>509.5,-86.5,509.5,-84</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>519.5,-86.5,519.5,-84</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>529.5,-86.5,529.5,-84</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>539.5,-86.5,539.5,-84</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>489.5,-86.5,489.5,-84</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>43</ID>
<points>477,-92.5,477.5,-92.5</points>
<connection>
<GID>747</GID>
<name>OUT</name></connection>
<intersection>477.5 27</intersection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-91.5,275.5,33</points>
<connection>
<GID>574</GID>
<name>OUT_0</name></connection>
<intersection>-91.5 16</intersection>
<intersection>-83.5 11</intersection>
<intersection>-59.5 3</intersection>
<intersection>-51.5 1</intersection>
<intersection>-17 34</intersection>
<intersection>-9 29</intersection>
<intersection>15 21</intersection>
<intersection>23 19</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-51.5,278.5,-51.5</points>
<connection>
<GID>575</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>275.5,-59.5,278.5,-59.5</points>
<connection>
<GID>612</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>275.5,-83.5,278.5,-83.5</points>
<connection>
<GID>699</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>275.5,-91.5,278.5,-91.5</points>
<connection>
<GID>746</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>275.5,23,278.5,23</points>
<connection>
<GID>556</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>275.5,15,278.5,15</points>
<connection>
<GID>558</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>275.5,-9,278.5,-9</points>
<connection>
<GID>564</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>275.5,-17,278.5,-17</points>
<connection>
<GID>566</GID>
<name>IN_2</name></connection>
<intersection>275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485.5,-97.5,485.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>485.5,-97.5,488.5,-97.5</points>
<intersection>485.5 0</intersection>
<intersection>488.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>485.5,-86.5,487.5,-86.5</points>
<connection>
<GID>743</GID>
<name>IN_1</name></connection>
<intersection>485.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>488.5,-100.5,488.5,-97.5</points>
<connection>
<GID>742</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>498.5,-92.5,499.5,-92.5</points>
<connection>
<GID>751</GID>
<name>IN_1</name></connection>
<connection>
<GID>749</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>501.5,-92.5,502.5,-92.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<connection>
<GID>750</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495.5,-97.5,495.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495.5,-97.5,498.5,-97.5</points>
<intersection>495.5 0</intersection>
<intersection>498.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>495.5,-86.5,497.5,-86.5</points>
<connection>
<GID>749</GID>
<name>IN_1</name></connection>
<intersection>495.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>498.5,-100.5,498.5,-97.5</points>
<connection>
<GID>748</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>508.5,-92.5,509.5,-92.5</points>
<connection>
<GID>755</GID>
<name>IN_1</name></connection>
<connection>
<GID>753</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>511.5,-92.5,512.5,-92.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<connection>
<GID>754</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>505.5,-97.5,505.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>505.5,-97.5,508.5,-97.5</points>
<intersection>505.5 0</intersection>
<intersection>508.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>505.5,-86.5,507.5,-86.5</points>
<connection>
<GID>753</GID>
<name>IN_1</name></connection>
<intersection>505.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>508.5,-100.5,508.5,-97.5</points>
<connection>
<GID>752</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>518.5,-92.5,519.5,-92.5</points>
<connection>
<GID>759</GID>
<name>IN_1</name></connection>
<connection>
<GID>757</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>521.5,-92.5,522.5,-92.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<connection>
<GID>758</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>515.5,-97.5,515.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>515.5,-97.5,518.5,-97.5</points>
<intersection>515.5 0</intersection>
<intersection>518.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>515.5,-86.5,517.5,-86.5</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<intersection>515.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>518.5,-100.5,518.5,-97.5</points>
<connection>
<GID>756</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>528.5,-92.5,529.5,-92.5</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<connection>
<GID>761</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>531.5,-92.5,532.5,-92.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<connection>
<GID>762</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>525.5,-97.5,525.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525.5,-97.5,528.5,-97.5</points>
<intersection>525.5 0</intersection>
<intersection>528.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525.5,-86.5,527.5,-86.5</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<intersection>525.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>528.5,-100.5,528.5,-97.5</points>
<connection>
<GID>760</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>538.5,-92.5,539.5,-92.5</points>
<connection>
<GID>767</GID>
<name>IN_1</name></connection>
<connection>
<GID>765</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>541.5,-92.5,542.5,-92.5</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<connection>
<GID>766</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535.5,-97.5,535.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535.5,-97.5,538.5,-97.5</points>
<intersection>535.5 0</intersection>
<intersection>538.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>535.5,-86.5,537.5,-86.5</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<intersection>535.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>538.5,-100.5,538.5,-97.5</points>
<connection>
<GID>764</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>548.5,-92.5,549.5,-92.5</points>
<connection>
<GID>771</GID>
<name>IN_1</name></connection>
<connection>
<GID>769</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>551.5,-92.5,552.5,-92.5</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<connection>
<GID>770</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>545.5,-97.5,545.5,-86.5</points>
<intersection>-97.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>545.5,-97.5,548.5,-97.5</points>
<intersection>545.5 0</intersection>
<intersection>548.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>545.5,-86.5,547.5,-86.5</points>
<connection>
<GID>769</GID>
<name>IN_1</name></connection>
<intersection>545.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>548.5,-100.5,548.5,-97.5</points>
<connection>
<GID>768</GID>
<name>OUT_0</name></connection>
<intersection>-97.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>482.5,-100.5,482.5,-83</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477,-83,482.5,-83</points>
<connection>
<GID>774</GID>
<name>OUT_0</name></connection>
<intersection>482.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,-73.5,273.5,33</points>
<connection>
<GID>572</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 7</intersection>
<intersection>-65.5 5</intersection>
<intersection>-57.5 3</intersection>
<intersection>-49.5 1</intersection>
<intersection>1 16</intersection>
<intersection>9 14</intersection>
<intersection>17 12</intersection>
<intersection>25 10</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273.5,-49.5,278.5,-49.5</points>
<connection>
<GID>575</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>273.5,-57.5,278.5,-57.5</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>273.5,-65.5,278.5,-65.5</points>
<connection>
<GID>630</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>273.5,-73.5,278.5,-73.5</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>273.5,25,278.5,25</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>273.5,17,278.5,17</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>273.5,9,278.5,9</points>
<connection>
<GID>560</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>273.5,1,278.5,1</points>
<connection>
<GID>562</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>490.5,-100.5,490.5,-98.5</points>
<connection>
<GID>745</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>490.5,-100.5,492.5,-100.5</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>490.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>742</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>510.5,-100.5,510.5,-98.5</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>510.5,-100.5,512.5,-100.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>510.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>500.5,-100.5,500.5,-98.5</points>
<connection>
<GID>751</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>500.5,-100.5,502.5,-100.5</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<intersection>500.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>744</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>520.5,-100.5,520.5,-98.5</points>
<connection>
<GID>759</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>520.5,-100.5,522.5,-100.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>520.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>745</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530.5,-100.5,530.5,-98.5</points>
<connection>
<GID>763</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530.5,-100.5,532.5,-100.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>530.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>746</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>540.5,-100.5,540.5,-98.5</points>
<connection>
<GID>767</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>540.5,-100.5,542.5,-100.5</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>540.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>747</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>550.5,-100.5,550.5,-98.5</points>
<connection>
<GID>771</GID>
<name>OUT</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>550.5,-100.5,552.5,-100.5</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<intersection>550.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>551.5,-86.5,551.5,-76</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-76,551.5,-76</points>
<connection>
<GID>774</GID>
<name>OUT_7</name></connection>
<intersection>551.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>749</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>541.5,-86.5,541.5,-77</points>
<connection>
<GID>766</GID>
<name>IN_1</name></connection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-77,541.5,-77</points>
<connection>
<GID>774</GID>
<name>OUT_6</name></connection>
<intersection>541.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>750</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531.5,-86.5,531.5,-78</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-78,531.5,-78</points>
<connection>
<GID>774</GID>
<name>OUT_5</name></connection>
<intersection>531.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>751</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>521.5,-86.5,521.5,-79</points>
<connection>
<GID>758</GID>
<name>IN_1</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-79,521.5,-79</points>
<connection>
<GID>774</GID>
<name>OUT_4</name></connection>
<intersection>521.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>752</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,-86.5,511.5,-80</points>
<connection>
<GID>754</GID>
<name>IN_1</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-80,511.5,-80</points>
<connection>
<GID>774</GID>
<name>OUT_3</name></connection>
<intersection>511.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>753</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501.5,-86.5,501.5,-81</points>
<connection>
<GID>750</GID>
<name>IN_1</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>477,-81,501.5,-81</points>
<connection>
<GID>774</GID>
<name>OUT_2</name></connection>
<intersection>501.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>754</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>472,-85,472,-85</points>
<connection>
<GID>774</GID>
<name>clock</name></connection>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>755</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,-86.5,468,-83</points>
<intersection>-86.5 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>468,-83,469,-83</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>468 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-86.5,468,-86.5</points>
<connection>
<GID>784</GID>
<name>OUT_0</name></connection>
<intersection>468 0</intersection></hsegment></shape></wire>
<wire>
<ID>756</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-84.5,467,-82</points>
<intersection>-84.5 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>464,-84.5,467,-84.5</points>
<connection>
<GID>783</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>467,-82,469,-82</points>
<connection>
<GID>774</GID>
<name>IN_1</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>757</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466,-82.5,466,-81</points>
<intersection>-82.5 2</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>466,-81,469,-81</points>
<connection>
<GID>774</GID>
<name>IN_2</name></connection>
<intersection>466 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-82.5,466,-82.5</points>
<connection>
<GID>782</GID>
<name>OUT_0</name></connection>
<intersection>466 0</intersection></hsegment></shape></wire>
<wire>
<ID>758</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,-80.5,465,-80</points>
<intersection>-80.5 3</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>465,-80,469,-80</points>
<connection>
<GID>774</GID>
<name>IN_3</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>464,-80.5,465,-80.5</points>
<connection>
<GID>781</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>759</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,-79,465,-78.5</points>
<intersection>-79 1</intersection>
<intersection>-78.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>465,-79,469,-79</points>
<connection>
<GID>774</GID>
<name>IN_4</name></connection>
<intersection>465 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>464,-78.5,465,-78.5</points>
<connection>
<GID>780</GID>
<name>OUT_0</name></connection>
<intersection>465 0</intersection></hsegment></shape></wire>
<wire>
<ID>760</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>467,-77,467,-74.5</points>
<intersection>-77 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467,-77,469,-77</points>
<connection>
<GID>774</GID>
<name>IN_6</name></connection>
<intersection>467 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>464,-74.5,467,-74.5</points>
<connection>
<GID>778</GID>
<name>OUT_0</name></connection>
<intersection>467 0</intersection></hsegment></shape></wire>
<wire>
<ID>761</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>466,-78,466,-76.5</points>
<intersection>-78 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>464,-76.5,466,-76.5</points>
<connection>
<GID>779</GID>
<name>OUT_0</name></connection>
<intersection>466 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>466,-78,469,-78</points>
<connection>
<GID>774</GID>
<name>IN_5</name></connection>
<intersection>466 0</intersection></hsegment></shape></wire>
<wire>
<ID>762</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>468,-76,468,-72.5</points>
<intersection>-76 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>464,-72.5,468,-72.5</points>
<connection>
<GID>777</GID>
<name>OUT_0</name></connection>
<intersection>468 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>468,-76,469,-76</points>
<connection>
<GID>774</GID>
<name>IN_7</name></connection>
<intersection>468 0</intersection></hsegment></shape></wire>
<wire>
<ID>763</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>472,-74,472,-74</points>
<connection>
<GID>774</GID>
<name>load</name></connection>
<connection>
<GID>776</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>764</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-71.5,571.5,-69.5</points>
<connection>
<GID>786</GID>
<name>IN_0</name></connection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>564.5,-71.5,571.5,-71.5</points>
<connection>
<GID>661</GID>
<name>OUT</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>765</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-63.5,571.5,-61.5</points>
<connection>
<GID>786</GID>
<name>OUT_0</name></connection>
<connection>
<GID>787</GID>
<name>IN_0</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>571.5,-62.5,582.5,-62.5</points>
<intersection>571.5 0</intersection>
<intersection>582.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>582.5,-62.5,582.5,-41.5</points>
<intersection>-62.5 1</intersection>
<intersection>-41.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>582.5,-41.5,583.5,-41.5</points>
<connection>
<GID>785</GID>
<name>IN_0</name></connection>
<intersection>582.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>766</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-55.5,571.5,-53.5</points>
<connection>
<GID>787</GID>
<name>OUT_0</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection>
<intersection>-54.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>571.5,-54.5,581.5,-54.5</points>
<intersection>571.5 0</intersection>
<intersection>581.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>581.5,-54.5,581.5,-40.5</points>
<intersection>-54.5 3</intersection>
<intersection>-40.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>581.5,-40.5,583.5,-40.5</points>
<connection>
<GID>785</GID>
<name>IN_1</name></connection>
<intersection>581.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>767</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-47.5,571.5,-45.5</points>
<connection>
<GID>788</GID>
<name>OUT_0</name></connection>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>-46.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>571.5,-46.5,580.5,-46.5</points>
<intersection>571.5 0</intersection>
<intersection>580.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>580.5,-46.5,580.5,-39.5</points>
<intersection>-46.5 6</intersection>
<intersection>-39.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>580.5,-39.5,583.5,-39.5</points>
<connection>
<GID>785</GID>
<name>IN_2</name></connection>
<intersection>580.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>768</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-39.5,571.5,-37.5</points>
<connection>
<GID>789</GID>
<name>OUT_0</name></connection>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>571.5,-38.5,583.5,-38.5</points>
<connection>
<GID>785</GID>
<name>IN_3</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 1>
<page 2>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 2>
<page 3>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 3>
<page 4>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 4>
<page 5>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 5>
<page 6>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 6>
<page 7>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 7>
<page 8>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 8>
<page 9>
<PageViewport>0,566.028,1778,-350.972</PageViewport></page 9></circuit>